//Teal 0x088 is the transparent color of sprite sheet.
module Background (
    input  logic clk, 
    input  logic [9:0] x, 
    input  logic [9:0] y, 
    output logic [11:0] out 
);
    assign logic[9:0] x_in = x;
    assign logic[9:0] y_in = y;
    assign logic[18:0] index = y_in * 640 + x_in;

always_ff @ (posedge clk)
    case (index)
      20'h00000: out <= 12'h222;
      20'h00001: out <= 12'h6af;
      20'h00002: out <= 12'h6af;
      20'h00003: out <= 12'h6af;
      20'h00004: out <= 12'h6af;
      20'h00005: out <= 12'h6af;
      20'h00006: out <= 12'h6af;
      20'h00007: out <= 12'h6af;
      20'h00008: out <= 12'h6af;
      20'h00009: out <= 12'h6af;
      20'h0000a: out <= 12'h6af;
      20'h0000b: out <= 12'h6af;
      20'h0000c: out <= 12'h6af;
      20'h0000d: out <= 12'h222;
      20'h0000e: out <= 12'h222;
      20'h0000f: out <= 12'h222;
      20'h00010: out <= 12'h000;
      20'h00011: out <= 12'h6af;
      20'h00012: out <= 12'h6af;
      20'h00013: out <= 12'h6af;
      20'h00014: out <= 12'h6af;
      20'h00015: out <= 12'h6af;
      20'h00016: out <= 12'h6af;
      20'h00017: out <= 12'h6af;
      20'h00018: out <= 12'h6af;
      20'h00019: out <= 12'h6af;
      20'h0001a: out <= 12'h6af;
      20'h0001b: out <= 12'h6af;
      20'h0001c: out <= 12'h6af;
      20'h0001d: out <= 12'h000;
      20'h0001e: out <= 12'h000;
      20'h0001f: out <= 12'h000;
      20'h00020: out <= 12'h222;
      20'h00021: out <= 12'h222;
      20'h00022: out <= 12'h222;
      20'h00023: out <= 12'h222;
      20'h00024: out <= 12'h222;
      20'h00025: out <= 12'h222;
      20'h00026: out <= 12'h222;
      20'h00027: out <= 12'h6af;
      20'h00028: out <= 12'hfff;
      20'h00029: out <= 12'h6af;
      20'h0002a: out <= 12'h222;
      20'h0002b: out <= 12'h222;
      20'h0002c: out <= 12'h222;
      20'h0002d: out <= 12'h222;
      20'h0002e: out <= 12'h222;
      20'h0002f: out <= 12'h222;
      20'h00030: out <= 12'h000;
      20'h00031: out <= 12'h000;
      20'h00032: out <= 12'h000;
      20'h00033: out <= 12'h000;
      20'h00034: out <= 12'h000;
      20'h00035: out <= 12'h000;
      20'h00036: out <= 12'h000;
      20'h00037: out <= 12'h6af;
      20'h00038: out <= 12'hfff;
      20'h00039: out <= 12'h6af;
      20'h0003a: out <= 12'h000;
      20'h0003b: out <= 12'h000;
      20'h0003c: out <= 12'h000;
      20'h0003d: out <= 12'h000;
      20'h0003e: out <= 12'h000;
      20'h0003f: out <= 12'h000;
      20'h00040: out <= 12'h222;
      20'h00041: out <= 12'h222;
      20'h00042: out <= 12'h222;
      20'h00043: out <= 12'h6af;
      20'h00044: out <= 12'h6af;
      20'h00045: out <= 12'h6af;
      20'h00046: out <= 12'h6af;
      20'h00047: out <= 12'h6af;
      20'h00048: out <= 12'h6af;
      20'h00049: out <= 12'h6af;
      20'h0004a: out <= 12'h6af;
      20'h0004b: out <= 12'h6af;
      20'h0004c: out <= 12'h6af;
      20'h0004d: out <= 12'h6af;
      20'h0004e: out <= 12'h6af;
      20'h0004f: out <= 12'h222;
      20'h00050: out <= 12'h000;
      20'h00051: out <= 12'h000;
      20'h00052: out <= 12'h000;
      20'h00053: out <= 12'h6af;
      20'h00054: out <= 12'h6af;
      20'h00055: out <= 12'h6af;
      20'h00056: out <= 12'h6af;
      20'h00057: out <= 12'h6af;
      20'h00058: out <= 12'h6af;
      20'h00059: out <= 12'h6af;
      20'h0005a: out <= 12'h6af;
      20'h0005b: out <= 12'h6af;
      20'h0005c: out <= 12'h6af;
      20'h0005d: out <= 12'h6af;
      20'h0005e: out <= 12'h6af;
      20'h0005f: out <= 12'h000;
      20'h00060: out <= 12'h222;
      20'h00061: out <= 12'h222;
      20'h00062: out <= 12'h222;
      20'h00063: out <= 12'h222;
      20'h00064: out <= 12'h222;
      20'h00065: out <= 12'h222;
      20'h00066: out <= 12'h222;
      20'h00067: out <= 12'h222;
      20'h00068: out <= 12'h222;
      20'h00069: out <= 12'h222;
      20'h0006a: out <= 12'h222;
      20'h0006b: out <= 12'h222;
      20'h0006c: out <= 12'h222;
      20'h0006d: out <= 12'h222;
      20'h0006e: out <= 12'h222;
      20'h0006f: out <= 12'h222;
      20'h00070: out <= 12'h000;
      20'h00071: out <= 12'h000;
      20'h00072: out <= 12'h000;
      20'h00073: out <= 12'h000;
      20'h00074: out <= 12'h000;
      20'h00075: out <= 12'h000;
      20'h00076: out <= 12'h000;
      20'h00077: out <= 12'h000;
      20'h00078: out <= 12'h000;
      20'h00079: out <= 12'h000;
      20'h0007a: out <= 12'h000;
      20'h0007b: out <= 12'h000;
      20'h0007c: out <= 12'h000;
      20'h0007d: out <= 12'h000;
      20'h0007e: out <= 12'h000;
      20'h0007f: out <= 12'h000;
      20'h00080: out <= 12'h603;
      20'h00081: out <= 12'h603;
      20'h00082: out <= 12'h603;
      20'h00083: out <= 12'h603;
      20'h00084: out <= 12'hee9;
      20'h00085: out <= 12'hee9;
      20'h00086: out <= 12'hee9;
      20'h00087: out <= 12'hee9;
      20'h00088: out <= 12'hb27;
      20'h00089: out <= 12'hee9;
      20'h0008a: out <= 12'hee9;
      20'h0008b: out <= 12'hee9;
      20'h0008c: out <= 12'hee9;
      20'h0008d: out <= 12'hee9;
      20'h0008e: out <= 12'hee9;
      20'h0008f: out <= 12'hee9;
      20'h00090: out <= 12'hb27;
      20'h00091: out <= 12'hee9;
      20'h00092: out <= 12'hee9;
      20'h00093: out <= 12'hee9;
      20'h00094: out <= 12'h000;
      20'h00095: out <= 12'h000;
      20'h00096: out <= 12'h000;
      20'h00097: out <= 12'h000;
      20'h00098: out <= 12'h000;
      20'h00099: out <= 12'h000;
      20'h0009a: out <= 12'h000;
      20'h0009b: out <= 12'h000;
      20'h0009c: out <= 12'hee9;
      20'h0009d: out <= 12'hee9;
      20'h0009e: out <= 12'hee9;
      20'h0009f: out <= 12'hee9;
      20'h000a0: out <= 12'hb27;
      20'h000a1: out <= 12'hee9;
      20'h000a2: out <= 12'hee9;
      20'h000a3: out <= 12'hee9;
      20'h000a4: out <= 12'h000;
      20'h000a5: out <= 12'h000;
      20'h000a6: out <= 12'h000;
      20'h000a7: out <= 12'h000;
      20'h000a8: out <= 12'h000;
      20'h000a9: out <= 12'h000;
      20'h000aa: out <= 12'h000;
      20'h000ab: out <= 12'h000;
      20'h000ac: out <= 12'h000;
      20'h000ad: out <= 12'h000;
      20'h000ae: out <= 12'h000;
      20'h000af: out <= 12'h000;
      20'h000b0: out <= 12'h000;
      20'h000b1: out <= 12'h000;
      20'h000b2: out <= 12'h000;
      20'h000b3: out <= 12'h000;
      20'h000b4: out <= 12'hee9;
      20'h000b5: out <= 12'hee9;
      20'h000b6: out <= 12'hee9;
      20'h000b7: out <= 12'hee9;
      20'h000b8: out <= 12'hb27;
      20'h000b9: out <= 12'hee9;
      20'h000ba: out <= 12'hee9;
      20'h000bb: out <= 12'hee9;
      20'h000bc: out <= 12'h000;
      20'h000bd: out <= 12'h000;
      20'h000be: out <= 12'h000;
      20'h000bf: out <= 12'h000;
      20'h000c0: out <= 12'h000;
      20'h000c1: out <= 12'h000;
      20'h000c2: out <= 12'h000;
      20'h000c3: out <= 12'h000;
      20'h000c4: out <= 12'hee9;
      20'h000c5: out <= 12'hee9;
      20'h000c6: out <= 12'hee9;
      20'h000c7: out <= 12'hee9;
      20'h000c8: out <= 12'hb27;
      20'h000c9: out <= 12'hee9;
      20'h000ca: out <= 12'hee9;
      20'h000cb: out <= 12'hee9;
      20'h000cc: out <= 12'hee9;
      20'h000cd: out <= 12'hee9;
      20'h000ce: out <= 12'hee9;
      20'h000cf: out <= 12'hee9;
      20'h000d0: out <= 12'hb27;
      20'h000d1: out <= 12'hee9;
      20'h000d2: out <= 12'hee9;
      20'h000d3: out <= 12'hee9;
      20'h000d4: out <= 12'h603;
      20'h000d5: out <= 12'h603;
      20'h000d6: out <= 12'h603;
      20'h000d7: out <= 12'h603;
      20'h000d8: out <= 12'hee9;
      20'h000d9: out <= 12'hee9;
      20'h000da: out <= 12'hee9;
      20'h000db: out <= 12'hee9;
      20'h000dc: out <= 12'hee9;
      20'h000dd: out <= 12'hee9;
      20'h000de: out <= 12'hee9;
      20'h000df: out <= 12'hb27;
      20'h000e0: out <= 12'hee9;
      20'h000e1: out <= 12'hee9;
      20'h000e2: out <= 12'hee9;
      20'h000e3: out <= 12'hee9;
      20'h000e4: out <= 12'hee9;
      20'h000e5: out <= 12'hee9;
      20'h000e6: out <= 12'hee9;
      20'h000e7: out <= 12'hb27;
      20'h000e8: out <= 12'hee9;
      20'h000e9: out <= 12'hee9;
      20'h000ea: out <= 12'hee9;
      20'h000eb: out <= 12'hee9;
      20'h000ec: out <= 12'hee9;
      20'h000ed: out <= 12'hee9;
      20'h000ee: out <= 12'hee9;
      20'h000ef: out <= 12'hb27;
      20'h000f0: out <= 12'hee9;
      20'h000f1: out <= 12'hee9;
      20'h000f2: out <= 12'hee9;
      20'h000f3: out <= 12'hee9;
      20'h000f4: out <= 12'hee9;
      20'h000f5: out <= 12'hee9;
      20'h000f6: out <= 12'hee9;
      20'h000f7: out <= 12'hb27;
      20'h000f8: out <= 12'hee9;
      20'h000f9: out <= 12'hee9;
      20'h000fa: out <= 12'hee9;
      20'h000fb: out <= 12'hee9;
      20'h000fc: out <= 12'hee9;
      20'h000fd: out <= 12'hee9;
      20'h000fe: out <= 12'hee9;
      20'h000ff: out <= 12'hb27;
      20'h00100: out <= 12'hee9;
      20'h00101: out <= 12'hee9;
      20'h00102: out <= 12'hee9;
      20'h00103: out <= 12'hee9;
      20'h00104: out <= 12'hee9;
      20'h00105: out <= 12'hee9;
      20'h00106: out <= 12'hee9;
      20'h00107: out <= 12'hb27;
      20'h00108: out <= 12'hee9;
      20'h00109: out <= 12'hee9;
      20'h0010a: out <= 12'hee9;
      20'h0010b: out <= 12'hee9;
      20'h0010c: out <= 12'hee9;
      20'h0010d: out <= 12'hee9;
      20'h0010e: out <= 12'hee9;
      20'h0010f: out <= 12'hb27;
      20'h00110: out <= 12'hee9;
      20'h00111: out <= 12'hee9;
      20'h00112: out <= 12'hee9;
      20'h00113: out <= 12'hee9;
      20'h00114: out <= 12'hee9;
      20'h00115: out <= 12'hee9;
      20'h00116: out <= 12'hee9;
      20'h00117: out <= 12'hb27;
      20'h00118: out <= 12'h222;
      20'h00119: out <= 12'hfff;
      20'h0011a: out <= 12'h16d;
      20'h0011b: out <= 12'hfff;
      20'h0011c: out <= 12'h16d;
      20'h0011d: out <= 12'hfff;
      20'h0011e: out <= 12'h16d;
      20'h0011f: out <= 12'hfff;
      20'h00120: out <= 12'h16d;
      20'h00121: out <= 12'hfff;
      20'h00122: out <= 12'h16d;
      20'h00123: out <= 12'hfff;
      20'h00124: out <= 12'h16d;
      20'h00125: out <= 12'h222;
      20'h00126: out <= 12'h222;
      20'h00127: out <= 12'h222;
      20'h00128: out <= 12'h000;
      20'h00129: out <= 12'h6af;
      20'h0012a: out <= 12'hfff;
      20'h0012b: out <= 12'h16d;
      20'h0012c: out <= 12'hfff;
      20'h0012d: out <= 12'h16d;
      20'h0012e: out <= 12'hfff;
      20'h0012f: out <= 12'h16d;
      20'h00130: out <= 12'hfff;
      20'h00131: out <= 12'h16d;
      20'h00132: out <= 12'hfff;
      20'h00133: out <= 12'h16d;
      20'h00134: out <= 12'hfff;
      20'h00135: out <= 12'h000;
      20'h00136: out <= 12'h000;
      20'h00137: out <= 12'h000;
      20'h00138: out <= 12'h222;
      20'h00139: out <= 12'h222;
      20'h0013a: out <= 12'h222;
      20'h0013b: out <= 12'h222;
      20'h0013c: out <= 12'h222;
      20'h0013d: out <= 12'h222;
      20'h0013e: out <= 12'h222;
      20'h0013f: out <= 12'h16d;
      20'h00140: out <= 12'hfff;
      20'h00141: out <= 12'h16d;
      20'h00142: out <= 12'h222;
      20'h00143: out <= 12'h222;
      20'h00144: out <= 12'h222;
      20'h00145: out <= 12'h222;
      20'h00146: out <= 12'h222;
      20'h00147: out <= 12'h222;
      20'h00148: out <= 12'h000;
      20'h00149: out <= 12'h000;
      20'h0014a: out <= 12'h000;
      20'h0014b: out <= 12'h000;
      20'h0014c: out <= 12'h000;
      20'h0014d: out <= 12'h000;
      20'h0014e: out <= 12'h000;
      20'h0014f: out <= 12'h16d;
      20'h00150: out <= 12'hfff;
      20'h00151: out <= 12'h16d;
      20'h00152: out <= 12'h000;
      20'h00153: out <= 12'h000;
      20'h00154: out <= 12'h000;
      20'h00155: out <= 12'h000;
      20'h00156: out <= 12'h000;
      20'h00157: out <= 12'h000;
      20'h00158: out <= 12'h222;
      20'h00159: out <= 12'h222;
      20'h0015a: out <= 12'h222;
      20'h0015b: out <= 12'h16d;
      20'h0015c: out <= 12'hfff;
      20'h0015d: out <= 12'h16d;
      20'h0015e: out <= 12'hfff;
      20'h0015f: out <= 12'h16d;
      20'h00160: out <= 12'hfff;
      20'h00161: out <= 12'h16d;
      20'h00162: out <= 12'hfff;
      20'h00163: out <= 12'h16d;
      20'h00164: out <= 12'hfff;
      20'h00165: out <= 12'h16d;
      20'h00166: out <= 12'hfff;
      20'h00167: out <= 12'h222;
      20'h00168: out <= 12'h000;
      20'h00169: out <= 12'h000;
      20'h0016a: out <= 12'h000;
      20'h0016b: out <= 12'hfff;
      20'h0016c: out <= 12'h16d;
      20'h0016d: out <= 12'hfff;
      20'h0016e: out <= 12'h16d;
      20'h0016f: out <= 12'hfff;
      20'h00170: out <= 12'h16d;
      20'h00171: out <= 12'hfff;
      20'h00172: out <= 12'h16d;
      20'h00173: out <= 12'hfff;
      20'h00174: out <= 12'h16d;
      20'h00175: out <= 12'hfff;
      20'h00176: out <= 12'h6af;
      20'h00177: out <= 12'h000;
      20'h00178: out <= 12'h222;
      20'h00179: out <= 12'h6af;
      20'h0017a: out <= 12'hfff;
      20'h0017b: out <= 12'h6af;
      20'h0017c: out <= 12'h222;
      20'h0017d: out <= 12'h222;
      20'h0017e: out <= 12'h222;
      20'h0017f: out <= 12'h222;
      20'h00180: out <= 12'h222;
      20'h00181: out <= 12'h222;
      20'h00182: out <= 12'h222;
      20'h00183: out <= 12'h222;
      20'h00184: out <= 12'h222;
      20'h00185: out <= 12'h6af;
      20'h00186: out <= 12'hfff;
      20'h00187: out <= 12'h6af;
      20'h00188: out <= 12'h000;
      20'h00189: out <= 12'h6af;
      20'h0018a: out <= 12'h6af;
      20'h0018b: out <= 12'h6af;
      20'h0018c: out <= 12'h000;
      20'h0018d: out <= 12'h000;
      20'h0018e: out <= 12'h000;
      20'h0018f: out <= 12'h000;
      20'h00190: out <= 12'h000;
      20'h00191: out <= 12'h000;
      20'h00192: out <= 12'h000;
      20'h00193: out <= 12'h000;
      20'h00194: out <= 12'h000;
      20'h00195: out <= 12'h6af;
      20'h00196: out <= 12'h6af;
      20'h00197: out <= 12'h6af;
      20'h00198: out <= 12'h603;
      20'h00199: out <= 12'h603;
      20'h0019a: out <= 12'h603;
      20'h0019b: out <= 12'h603;
      20'h0019c: out <= 12'hf87;
      20'h0019d: out <= 12'hf87;
      20'h0019e: out <= 12'hf87;
      20'h0019f: out <= 12'hee9;
      20'h001a0: out <= 12'hb27;
      20'h001a1: out <= 12'hf87;
      20'h001a2: out <= 12'hf87;
      20'h001a3: out <= 12'hf87;
      20'h001a4: out <= 12'hf87;
      20'h001a5: out <= 12'hf87;
      20'h001a6: out <= 12'hf87;
      20'h001a7: out <= 12'hee9;
      20'h001a8: out <= 12'hb27;
      20'h001a9: out <= 12'hf87;
      20'h001aa: out <= 12'hf87;
      20'h001ab: out <= 12'hf87;
      20'h001ac: out <= 12'h000;
      20'h001ad: out <= 12'h000;
      20'h001ae: out <= 12'h000;
      20'h001af: out <= 12'h000;
      20'h001b0: out <= 12'h000;
      20'h001b1: out <= 12'h000;
      20'h001b2: out <= 12'h000;
      20'h001b3: out <= 12'h000;
      20'h001b4: out <= 12'hf87;
      20'h001b5: out <= 12'hf87;
      20'h001b6: out <= 12'hf87;
      20'h001b7: out <= 12'hee9;
      20'h001b8: out <= 12'hb27;
      20'h001b9: out <= 12'hf87;
      20'h001ba: out <= 12'hf87;
      20'h001bb: out <= 12'hf87;
      20'h001bc: out <= 12'h000;
      20'h001bd: out <= 12'h000;
      20'h001be: out <= 12'h000;
      20'h001bf: out <= 12'h000;
      20'h001c0: out <= 12'h000;
      20'h001c1: out <= 12'h000;
      20'h001c2: out <= 12'h000;
      20'h001c3: out <= 12'h000;
      20'h001c4: out <= 12'h000;
      20'h001c5: out <= 12'h000;
      20'h001c6: out <= 12'h000;
      20'h001c7: out <= 12'h000;
      20'h001c8: out <= 12'h000;
      20'h001c9: out <= 12'h000;
      20'h001ca: out <= 12'h000;
      20'h001cb: out <= 12'h000;
      20'h001cc: out <= 12'hf87;
      20'h001cd: out <= 12'hf87;
      20'h001ce: out <= 12'hf87;
      20'h001cf: out <= 12'hee9;
      20'h001d0: out <= 12'hb27;
      20'h001d1: out <= 12'hf87;
      20'h001d2: out <= 12'hf87;
      20'h001d3: out <= 12'hf87;
      20'h001d4: out <= 12'h000;
      20'h001d5: out <= 12'h000;
      20'h001d6: out <= 12'h000;
      20'h001d7: out <= 12'h000;
      20'h001d8: out <= 12'h000;
      20'h001d9: out <= 12'h000;
      20'h001da: out <= 12'h000;
      20'h001db: out <= 12'h000;
      20'h001dc: out <= 12'hf87;
      20'h001dd: out <= 12'hf87;
      20'h001de: out <= 12'hf87;
      20'h001df: out <= 12'hee9;
      20'h001e0: out <= 12'hb27;
      20'h001e1: out <= 12'hf87;
      20'h001e2: out <= 12'hf87;
      20'h001e3: out <= 12'hf87;
      20'h001e4: out <= 12'hf87;
      20'h001e5: out <= 12'hf87;
      20'h001e6: out <= 12'hf87;
      20'h001e7: out <= 12'hee9;
      20'h001e8: out <= 12'hb27;
      20'h001e9: out <= 12'hf87;
      20'h001ea: out <= 12'hf87;
      20'h001eb: out <= 12'hf87;
      20'h001ec: out <= 12'h603;
      20'h001ed: out <= 12'h603;
      20'h001ee: out <= 12'h603;
      20'h001ef: out <= 12'h603;
      20'h001f0: out <= 12'hee9;
      20'h001f1: out <= 12'hf87;
      20'h001f2: out <= 12'hf87;
      20'h001f3: out <= 12'hf87;
      20'h001f4: out <= 12'hf87;
      20'h001f5: out <= 12'hf87;
      20'h001f6: out <= 12'hf87;
      20'h001f7: out <= 12'hb27;
      20'h001f8: out <= 12'hee9;
      20'h001f9: out <= 12'hf87;
      20'h001fa: out <= 12'hf87;
      20'h001fb: out <= 12'hf87;
      20'h001fc: out <= 12'hf87;
      20'h001fd: out <= 12'hf87;
      20'h001fe: out <= 12'hf87;
      20'h001ff: out <= 12'hb27;
      20'h00200: out <= 12'hee9;
      20'h00201: out <= 12'hf87;
      20'h00202: out <= 12'hf87;
      20'h00203: out <= 12'hf87;
      20'h00204: out <= 12'hf87;
      20'h00205: out <= 12'hf87;
      20'h00206: out <= 12'hf87;
      20'h00207: out <= 12'hb27;
      20'h00208: out <= 12'hee9;
      20'h00209: out <= 12'hf87;
      20'h0020a: out <= 12'hf87;
      20'h0020b: out <= 12'hf87;
      20'h0020c: out <= 12'hf87;
      20'h0020d: out <= 12'hf87;
      20'h0020e: out <= 12'hf87;
      20'h0020f: out <= 12'hb27;
      20'h00210: out <= 12'hee9;
      20'h00211: out <= 12'hf87;
      20'h00212: out <= 12'hf87;
      20'h00213: out <= 12'hf87;
      20'h00214: out <= 12'hf87;
      20'h00215: out <= 12'hf87;
      20'h00216: out <= 12'hf87;
      20'h00217: out <= 12'hb27;
      20'h00218: out <= 12'hee9;
      20'h00219: out <= 12'hf87;
      20'h0021a: out <= 12'hf87;
      20'h0021b: out <= 12'hf87;
      20'h0021c: out <= 12'hf87;
      20'h0021d: out <= 12'hf87;
      20'h0021e: out <= 12'hf87;
      20'h0021f: out <= 12'hb27;
      20'h00220: out <= 12'hee9;
      20'h00221: out <= 12'hf87;
      20'h00222: out <= 12'hf87;
      20'h00223: out <= 12'hf87;
      20'h00224: out <= 12'hf87;
      20'h00225: out <= 12'hf87;
      20'h00226: out <= 12'hf87;
      20'h00227: out <= 12'hb27;
      20'h00228: out <= 12'hee9;
      20'h00229: out <= 12'hf87;
      20'h0022a: out <= 12'hf87;
      20'h0022b: out <= 12'hf87;
      20'h0022c: out <= 12'hf87;
      20'h0022d: out <= 12'hf87;
      20'h0022e: out <= 12'hf87;
      20'h0022f: out <= 12'hb27;
      20'h00230: out <= 12'h222;
      20'h00231: out <= 12'h6af;
      20'h00232: out <= 12'h6af;
      20'h00233: out <= 12'h6af;
      20'h00234: out <= 12'h16d;
      20'h00235: out <= 12'h16d;
      20'h00236: out <= 12'h16d;
      20'h00237: out <= 12'h16d;
      20'h00238: out <= 12'h16d;
      20'h00239: out <= 12'h16d;
      20'h0023a: out <= 12'h16d;
      20'h0023b: out <= 12'h6af;
      20'h0023c: out <= 12'h6af;
      20'h0023d: out <= 12'h222;
      20'h0023e: out <= 12'h222;
      20'h0023f: out <= 12'h222;
      20'h00240: out <= 12'h000;
      20'h00241: out <= 12'h6af;
      20'h00242: out <= 12'h6af;
      20'h00243: out <= 12'h6af;
      20'h00244: out <= 12'h16d;
      20'h00245: out <= 12'h16d;
      20'h00246: out <= 12'h16d;
      20'h00247: out <= 12'h16d;
      20'h00248: out <= 12'h16d;
      20'h00249: out <= 12'h16d;
      20'h0024a: out <= 12'h16d;
      20'h0024b: out <= 12'h6af;
      20'h0024c: out <= 12'h6af;
      20'h0024d: out <= 12'h000;
      20'h0024e: out <= 12'h000;
      20'h0024f: out <= 12'h000;
      20'h00250: out <= 12'h222;
      20'h00251: out <= 12'h222;
      20'h00252: out <= 12'h222;
      20'h00253: out <= 12'h222;
      20'h00254: out <= 12'h222;
      20'h00255: out <= 12'h222;
      20'h00256: out <= 12'h222;
      20'h00257: out <= 12'h16d;
      20'h00258: out <= 12'hfff;
      20'h00259: out <= 12'h16d;
      20'h0025a: out <= 12'h222;
      20'h0025b: out <= 12'h222;
      20'h0025c: out <= 12'h222;
      20'h0025d: out <= 12'h222;
      20'h0025e: out <= 12'h222;
      20'h0025f: out <= 12'h222;
      20'h00260: out <= 12'h000;
      20'h00261: out <= 12'h000;
      20'h00262: out <= 12'h000;
      20'h00263: out <= 12'h000;
      20'h00264: out <= 12'h000;
      20'h00265: out <= 12'h000;
      20'h00266: out <= 12'h000;
      20'h00267: out <= 12'h16d;
      20'h00268: out <= 12'hfff;
      20'h00269: out <= 12'h16d;
      20'h0026a: out <= 12'h000;
      20'h0026b: out <= 12'h000;
      20'h0026c: out <= 12'h000;
      20'h0026d: out <= 12'h000;
      20'h0026e: out <= 12'h000;
      20'h0026f: out <= 12'h000;
      20'h00270: out <= 12'h222;
      20'h00271: out <= 12'h222;
      20'h00272: out <= 12'h222;
      20'h00273: out <= 12'h6af;
      20'h00274: out <= 12'h6af;
      20'h00275: out <= 12'h16d;
      20'h00276: out <= 12'h16d;
      20'h00277: out <= 12'h16d;
      20'h00278: out <= 12'h16d;
      20'h00279: out <= 12'h16d;
      20'h0027a: out <= 12'h16d;
      20'h0027b: out <= 12'h16d;
      20'h0027c: out <= 12'h6af;
      20'h0027d: out <= 12'h6af;
      20'h0027e: out <= 12'h6af;
      20'h0027f: out <= 12'h222;
      20'h00280: out <= 12'h000;
      20'h00281: out <= 12'h000;
      20'h00282: out <= 12'h000;
      20'h00283: out <= 12'h6af;
      20'h00284: out <= 12'h6af;
      20'h00285: out <= 12'h16d;
      20'h00286: out <= 12'h16d;
      20'h00287: out <= 12'h16d;
      20'h00288: out <= 12'h16d;
      20'h00289: out <= 12'h16d;
      20'h0028a: out <= 12'h16d;
      20'h0028b: out <= 12'h16d;
      20'h0028c: out <= 12'h6af;
      20'h0028d: out <= 12'h6af;
      20'h0028e: out <= 12'h6af;
      20'h0028f: out <= 12'h000;
      20'h00290: out <= 12'h222;
      20'h00291: out <= 12'h6af;
      20'h00292: out <= 12'h16d;
      20'h00293: out <= 12'h6af;
      20'h00294: out <= 12'h222;
      20'h00295: out <= 12'h16d;
      20'h00296: out <= 12'h16d;
      20'h00297: out <= 12'h16d;
      20'h00298: out <= 12'h16d;
      20'h00299: out <= 12'h16d;
      20'h0029a: out <= 12'h16d;
      20'h0029b: out <= 12'h16d;
      20'h0029c: out <= 12'h222;
      20'h0029d: out <= 12'h6af;
      20'h0029e: out <= 12'h16d;
      20'h0029f: out <= 12'h6af;
      20'h002a0: out <= 12'h000;
      20'h002a1: out <= 12'h6af;
      20'h002a2: out <= 12'hfff;
      20'h002a3: out <= 12'h6af;
      20'h002a4: out <= 12'h000;
      20'h002a5: out <= 12'h16d;
      20'h002a6: out <= 12'h16d;
      20'h002a7: out <= 12'h16d;
      20'h002a8: out <= 12'h16d;
      20'h002a9: out <= 12'h16d;
      20'h002aa: out <= 12'h16d;
      20'h002ab: out <= 12'h16d;
      20'h002ac: out <= 12'h000;
      20'h002ad: out <= 12'h6af;
      20'h002ae: out <= 12'hfff;
      20'h002af: out <= 12'h6af;
      20'h002b0: out <= 12'h603;
      20'h002b1: out <= 12'h603;
      20'h002b2: out <= 12'h603;
      20'h002b3: out <= 12'h603;
      20'h002b4: out <= 12'hf87;
      20'h002b5: out <= 12'hf87;
      20'h002b6: out <= 12'hf87;
      20'h002b7: out <= 12'hee9;
      20'h002b8: out <= 12'hb27;
      20'h002b9: out <= 12'hf87;
      20'h002ba: out <= 12'hf87;
      20'h002bb: out <= 12'hf87;
      20'h002bc: out <= 12'hf87;
      20'h002bd: out <= 12'hf87;
      20'h002be: out <= 12'hf87;
      20'h002bf: out <= 12'hee9;
      20'h002c0: out <= 12'hb27;
      20'h002c1: out <= 12'hf87;
      20'h002c2: out <= 12'hf87;
      20'h002c3: out <= 12'hf87;
      20'h002c4: out <= 12'h000;
      20'h002c5: out <= 12'h000;
      20'h002c6: out <= 12'h000;
      20'h002c7: out <= 12'h000;
      20'h002c8: out <= 12'h000;
      20'h002c9: out <= 12'h000;
      20'h002ca: out <= 12'h000;
      20'h002cb: out <= 12'h000;
      20'h002cc: out <= 12'hf87;
      20'h002cd: out <= 12'hf87;
      20'h002ce: out <= 12'hf87;
      20'h002cf: out <= 12'hee9;
      20'h002d0: out <= 12'hb27;
      20'h002d1: out <= 12'hf87;
      20'h002d2: out <= 12'hf87;
      20'h002d3: out <= 12'hf87;
      20'h002d4: out <= 12'h000;
      20'h002d5: out <= 12'h000;
      20'h002d6: out <= 12'h000;
      20'h002d7: out <= 12'h000;
      20'h002d8: out <= 12'h000;
      20'h002d9: out <= 12'h000;
      20'h002da: out <= 12'h000;
      20'h002db: out <= 12'h000;
      20'h002dc: out <= 12'h000;
      20'h002dd: out <= 12'h000;
      20'h002de: out <= 12'h000;
      20'h002df: out <= 12'h000;
      20'h002e0: out <= 12'h000;
      20'h002e1: out <= 12'h000;
      20'h002e2: out <= 12'h000;
      20'h002e3: out <= 12'h000;
      20'h002e4: out <= 12'hf87;
      20'h002e5: out <= 12'hf87;
      20'h002e6: out <= 12'hf87;
      20'h002e7: out <= 12'hee9;
      20'h002e8: out <= 12'hb27;
      20'h002e9: out <= 12'hf87;
      20'h002ea: out <= 12'hf87;
      20'h002eb: out <= 12'hf87;
      20'h002ec: out <= 12'h000;
      20'h002ed: out <= 12'h000;
      20'h002ee: out <= 12'h000;
      20'h002ef: out <= 12'h000;
      20'h002f0: out <= 12'h000;
      20'h002f1: out <= 12'h000;
      20'h002f2: out <= 12'h000;
      20'h002f3: out <= 12'h000;
      20'h002f4: out <= 12'hf87;
      20'h002f5: out <= 12'hf87;
      20'h002f6: out <= 12'hf87;
      20'h002f7: out <= 12'hee9;
      20'h002f8: out <= 12'hb27;
      20'h002f9: out <= 12'hf87;
      20'h002fa: out <= 12'hf87;
      20'h002fb: out <= 12'hf87;
      20'h002fc: out <= 12'hf87;
      20'h002fd: out <= 12'hf87;
      20'h002fe: out <= 12'hf87;
      20'h002ff: out <= 12'hee9;
      20'h00300: out <= 12'hb27;
      20'h00301: out <= 12'hf87;
      20'h00302: out <= 12'hf87;
      20'h00303: out <= 12'hf87;
      20'h00304: out <= 12'h603;
      20'h00305: out <= 12'h603;
      20'h00306: out <= 12'h603;
      20'h00307: out <= 12'h603;
      20'h00308: out <= 12'hee9;
      20'h00309: out <= 12'hf87;
      20'h0030a: out <= 12'hee9;
      20'h0030b: out <= 12'hee9;
      20'h0030c: out <= 12'hee9;
      20'h0030d: out <= 12'hb27;
      20'h0030e: out <= 12'hf87;
      20'h0030f: out <= 12'hb27;
      20'h00310: out <= 12'hee9;
      20'h00311: out <= 12'hf87;
      20'h00312: out <= 12'hee9;
      20'h00313: out <= 12'hee9;
      20'h00314: out <= 12'hee9;
      20'h00315: out <= 12'hb27;
      20'h00316: out <= 12'hf87;
      20'h00317: out <= 12'hb27;
      20'h00318: out <= 12'hee9;
      20'h00319: out <= 12'hf87;
      20'h0031a: out <= 12'hee9;
      20'h0031b: out <= 12'hee9;
      20'h0031c: out <= 12'hee9;
      20'h0031d: out <= 12'hb27;
      20'h0031e: out <= 12'hf87;
      20'h0031f: out <= 12'hb27;
      20'h00320: out <= 12'hee9;
      20'h00321: out <= 12'hf87;
      20'h00322: out <= 12'hee9;
      20'h00323: out <= 12'hee9;
      20'h00324: out <= 12'hee9;
      20'h00325: out <= 12'hb27;
      20'h00326: out <= 12'hf87;
      20'h00327: out <= 12'hb27;
      20'h00328: out <= 12'hee9;
      20'h00329: out <= 12'hf87;
      20'h0032a: out <= 12'hee9;
      20'h0032b: out <= 12'hee9;
      20'h0032c: out <= 12'hee9;
      20'h0032d: out <= 12'hb27;
      20'h0032e: out <= 12'hf87;
      20'h0032f: out <= 12'hb27;
      20'h00330: out <= 12'hee9;
      20'h00331: out <= 12'hf87;
      20'h00332: out <= 12'hee9;
      20'h00333: out <= 12'hee9;
      20'h00334: out <= 12'hee9;
      20'h00335: out <= 12'hb27;
      20'h00336: out <= 12'hf87;
      20'h00337: out <= 12'hb27;
      20'h00338: out <= 12'hee9;
      20'h00339: out <= 12'hf87;
      20'h0033a: out <= 12'hee9;
      20'h0033b: out <= 12'hee9;
      20'h0033c: out <= 12'hee9;
      20'h0033d: out <= 12'hb27;
      20'h0033e: out <= 12'hf87;
      20'h0033f: out <= 12'hb27;
      20'h00340: out <= 12'hee9;
      20'h00341: out <= 12'hf87;
      20'h00342: out <= 12'hee9;
      20'h00343: out <= 12'hee9;
      20'h00344: out <= 12'hee9;
      20'h00345: out <= 12'hb27;
      20'h00346: out <= 12'hf87;
      20'h00347: out <= 12'hb27;
      20'h00348: out <= 12'h222;
      20'h00349: out <= 12'h222;
      20'h0034a: out <= 12'h222;
      20'h0034b: out <= 12'h16d;
      20'h0034c: out <= 12'hfff;
      20'h0034d: out <= 12'h6af;
      20'h0034e: out <= 12'h6af;
      20'h0034f: out <= 12'h6af;
      20'h00350: out <= 12'h6af;
      20'h00351: out <= 12'hfff;
      20'h00352: out <= 12'h16d;
      20'h00353: out <= 12'h222;
      20'h00354: out <= 12'h222;
      20'h00355: out <= 12'h222;
      20'h00356: out <= 12'h222;
      20'h00357: out <= 12'h222;
      20'h00358: out <= 12'h000;
      20'h00359: out <= 12'h000;
      20'h0035a: out <= 12'h000;
      20'h0035b: out <= 12'h16d;
      20'h0035c: out <= 12'hfff;
      20'h0035d: out <= 12'h6af;
      20'h0035e: out <= 12'h6af;
      20'h0035f: out <= 12'h6af;
      20'h00360: out <= 12'h6af;
      20'h00361: out <= 12'hfff;
      20'h00362: out <= 12'h16d;
      20'h00363: out <= 12'h000;
      20'h00364: out <= 12'h000;
      20'h00365: out <= 12'h000;
      20'h00366: out <= 12'h000;
      20'h00367: out <= 12'h000;
      20'h00368: out <= 12'h222;
      20'h00369: out <= 12'h6af;
      20'h0036a: out <= 12'h16d;
      20'h0036b: out <= 12'h6af;
      20'h0036c: out <= 12'h222;
      20'h0036d: out <= 12'h222;
      20'h0036e: out <= 12'h222;
      20'h0036f: out <= 12'h16d;
      20'h00370: out <= 12'hfff;
      20'h00371: out <= 12'h16d;
      20'h00372: out <= 12'h222;
      20'h00373: out <= 12'h222;
      20'h00374: out <= 12'h222;
      20'h00375: out <= 12'h6af;
      20'h00376: out <= 12'h16d;
      20'h00377: out <= 12'h6af;
      20'h00378: out <= 12'h000;
      20'h00379: out <= 12'h6af;
      20'h0037a: out <= 12'hfff;
      20'h0037b: out <= 12'h6af;
      20'h0037c: out <= 12'h000;
      20'h0037d: out <= 12'h000;
      20'h0037e: out <= 12'h000;
      20'h0037f: out <= 12'h16d;
      20'h00380: out <= 12'hfff;
      20'h00381: out <= 12'h16d;
      20'h00382: out <= 12'h000;
      20'h00383: out <= 12'h000;
      20'h00384: out <= 12'h000;
      20'h00385: out <= 12'h6af;
      20'h00386: out <= 12'hfff;
      20'h00387: out <= 12'h6af;
      20'h00388: out <= 12'h222;
      20'h00389: out <= 12'h222;
      20'h0038a: out <= 12'h222;
      20'h0038b: out <= 12'h222;
      20'h0038c: out <= 12'h222;
      20'h0038d: out <= 12'h16d;
      20'h0038e: out <= 12'hfff;
      20'h0038f: out <= 12'h6af;
      20'h00390: out <= 12'h6af;
      20'h00391: out <= 12'h6af;
      20'h00392: out <= 12'h6af;
      20'h00393: out <= 12'hfff;
      20'h00394: out <= 12'h16d;
      20'h00395: out <= 12'h222;
      20'h00396: out <= 12'h222;
      20'h00397: out <= 12'h222;
      20'h00398: out <= 12'h000;
      20'h00399: out <= 12'h000;
      20'h0039a: out <= 12'h000;
      20'h0039b: out <= 12'h000;
      20'h0039c: out <= 12'h000;
      20'h0039d: out <= 12'h16d;
      20'h0039e: out <= 12'hfff;
      20'h0039f: out <= 12'h6af;
      20'h003a0: out <= 12'h6af;
      20'h003a1: out <= 12'h6af;
      20'h003a2: out <= 12'h6af;
      20'h003a3: out <= 12'hfff;
      20'h003a4: out <= 12'h16d;
      20'h003a5: out <= 12'h000;
      20'h003a6: out <= 12'h000;
      20'h003a7: out <= 12'h000;
      20'h003a8: out <= 12'h222;
      20'h003a9: out <= 12'h6af;
      20'h003aa: out <= 12'hfff;
      20'h003ab: out <= 12'h6af;
      20'h003ac: out <= 12'h16d;
      20'h003ad: out <= 12'hfff;
      20'h003ae: out <= 12'h6af;
      20'h003af: out <= 12'h6af;
      20'h003b0: out <= 12'h6af;
      20'h003b1: out <= 12'h6af;
      20'h003b2: out <= 12'h6af;
      20'h003b3: out <= 12'hfff;
      20'h003b4: out <= 12'h16d;
      20'h003b5: out <= 12'h6af;
      20'h003b6: out <= 12'hfff;
      20'h003b7: out <= 12'h6af;
      20'h003b8: out <= 12'h000;
      20'h003b9: out <= 12'h6af;
      20'h003ba: out <= 12'h16d;
      20'h003bb: out <= 12'h6af;
      20'h003bc: out <= 12'h16d;
      20'h003bd: out <= 12'hfff;
      20'h003be: out <= 12'h6af;
      20'h003bf: out <= 12'h6af;
      20'h003c0: out <= 12'h6af;
      20'h003c1: out <= 12'h6af;
      20'h003c2: out <= 12'h6af;
      20'h003c3: out <= 12'hfff;
      20'h003c4: out <= 12'h16d;
      20'h003c5: out <= 12'h6af;
      20'h003c6: out <= 12'h16d;
      20'h003c7: out <= 12'h6af;
      20'h003c8: out <= 12'h603;
      20'h003c9: out <= 12'h603;
      20'h003ca: out <= 12'h603;
      20'h003cb: out <= 12'h603;
      20'h003cc: out <= 12'hb27;
      20'h003cd: out <= 12'hb27;
      20'h003ce: out <= 12'hb27;
      20'h003cf: out <= 12'hb27;
      20'h003d0: out <= 12'hb27;
      20'h003d1: out <= 12'hb27;
      20'h003d2: out <= 12'hb27;
      20'h003d3: out <= 12'hb27;
      20'h003d4: out <= 12'hb27;
      20'h003d5: out <= 12'hb27;
      20'h003d6: out <= 12'hb27;
      20'h003d7: out <= 12'hb27;
      20'h003d8: out <= 12'hb27;
      20'h003d9: out <= 12'hb27;
      20'h003da: out <= 12'hb27;
      20'h003db: out <= 12'hb27;
      20'h003dc: out <= 12'h000;
      20'h003dd: out <= 12'h000;
      20'h003de: out <= 12'h000;
      20'h003df: out <= 12'h000;
      20'h003e0: out <= 12'h000;
      20'h003e1: out <= 12'h000;
      20'h003e2: out <= 12'h000;
      20'h003e3: out <= 12'h000;
      20'h003e4: out <= 12'hb27;
      20'h003e5: out <= 12'hb27;
      20'h003e6: out <= 12'hb27;
      20'h003e7: out <= 12'hb27;
      20'h003e8: out <= 12'hb27;
      20'h003e9: out <= 12'hb27;
      20'h003ea: out <= 12'hb27;
      20'h003eb: out <= 12'hb27;
      20'h003ec: out <= 12'h000;
      20'h003ed: out <= 12'h000;
      20'h003ee: out <= 12'h000;
      20'h003ef: out <= 12'h000;
      20'h003f0: out <= 12'h000;
      20'h003f1: out <= 12'h000;
      20'h003f2: out <= 12'h000;
      20'h003f3: out <= 12'h000;
      20'h003f4: out <= 12'h000;
      20'h003f5: out <= 12'h000;
      20'h003f6: out <= 12'h000;
      20'h003f7: out <= 12'h000;
      20'h003f8: out <= 12'h000;
      20'h003f9: out <= 12'h000;
      20'h003fa: out <= 12'h000;
      20'h003fb: out <= 12'h000;
      20'h003fc: out <= 12'hb27;
      20'h003fd: out <= 12'hb27;
      20'h003fe: out <= 12'hb27;
      20'h003ff: out <= 12'hb27;
      20'h00400: out <= 12'hb27;
      20'h00401: out <= 12'hb27;
      20'h00402: out <= 12'hb27;
      20'h00403: out <= 12'hb27;
      20'h00404: out <= 12'h000;
      20'h00405: out <= 12'h000;
      20'h00406: out <= 12'h000;
      20'h00407: out <= 12'h000;
      20'h00408: out <= 12'h000;
      20'h00409: out <= 12'h000;
      20'h0040a: out <= 12'h000;
      20'h0040b: out <= 12'h000;
      20'h0040c: out <= 12'hb27;
      20'h0040d: out <= 12'hb27;
      20'h0040e: out <= 12'hb27;
      20'h0040f: out <= 12'hb27;
      20'h00410: out <= 12'hb27;
      20'h00411: out <= 12'hb27;
      20'h00412: out <= 12'hb27;
      20'h00413: out <= 12'hb27;
      20'h00414: out <= 12'hb27;
      20'h00415: out <= 12'hb27;
      20'h00416: out <= 12'hb27;
      20'h00417: out <= 12'hb27;
      20'h00418: out <= 12'hb27;
      20'h00419: out <= 12'hb27;
      20'h0041a: out <= 12'hb27;
      20'h0041b: out <= 12'hb27;
      20'h0041c: out <= 12'h603;
      20'h0041d: out <= 12'h603;
      20'h0041e: out <= 12'h603;
      20'h0041f: out <= 12'h603;
      20'h00420: out <= 12'hee9;
      20'h00421: out <= 12'hf87;
      20'h00422: out <= 12'hee9;
      20'h00423: out <= 12'hf87;
      20'h00424: out <= 12'hf87;
      20'h00425: out <= 12'hb27;
      20'h00426: out <= 12'hf87;
      20'h00427: out <= 12'hb27;
      20'h00428: out <= 12'hee9;
      20'h00429: out <= 12'hf87;
      20'h0042a: out <= 12'hee9;
      20'h0042b: out <= 12'hf87;
      20'h0042c: out <= 12'hf87;
      20'h0042d: out <= 12'hb27;
      20'h0042e: out <= 12'hf87;
      20'h0042f: out <= 12'hb27;
      20'h00430: out <= 12'hee9;
      20'h00431: out <= 12'hf87;
      20'h00432: out <= 12'hee9;
      20'h00433: out <= 12'hf87;
      20'h00434: out <= 12'hf87;
      20'h00435: out <= 12'hb27;
      20'h00436: out <= 12'hf87;
      20'h00437: out <= 12'hb27;
      20'h00438: out <= 12'hee9;
      20'h00439: out <= 12'hf87;
      20'h0043a: out <= 12'hee9;
      20'h0043b: out <= 12'hf87;
      20'h0043c: out <= 12'hf87;
      20'h0043d: out <= 12'hb27;
      20'h0043e: out <= 12'hf87;
      20'h0043f: out <= 12'hb27;
      20'h00440: out <= 12'hee9;
      20'h00441: out <= 12'hf87;
      20'h00442: out <= 12'hee9;
      20'h00443: out <= 12'hf87;
      20'h00444: out <= 12'hf87;
      20'h00445: out <= 12'hb27;
      20'h00446: out <= 12'hf87;
      20'h00447: out <= 12'hb27;
      20'h00448: out <= 12'hee9;
      20'h00449: out <= 12'hf87;
      20'h0044a: out <= 12'hee9;
      20'h0044b: out <= 12'hf87;
      20'h0044c: out <= 12'hf87;
      20'h0044d: out <= 12'hb27;
      20'h0044e: out <= 12'hf87;
      20'h0044f: out <= 12'hb27;
      20'h00450: out <= 12'hee9;
      20'h00451: out <= 12'hf87;
      20'h00452: out <= 12'hee9;
      20'h00453: out <= 12'hf87;
      20'h00454: out <= 12'hf87;
      20'h00455: out <= 12'hb27;
      20'h00456: out <= 12'hf87;
      20'h00457: out <= 12'hb27;
      20'h00458: out <= 12'hee9;
      20'h00459: out <= 12'hf87;
      20'h0045a: out <= 12'hee9;
      20'h0045b: out <= 12'hf87;
      20'h0045c: out <= 12'hf87;
      20'h0045d: out <= 12'hb27;
      20'h0045e: out <= 12'hf87;
      20'h0045f: out <= 12'hb27;
      20'h00460: out <= 12'h222;
      20'h00461: out <= 12'h222;
      20'h00462: out <= 12'h16d;
      20'h00463: out <= 12'hfff;
      20'h00464: out <= 12'h6af;
      20'h00465: out <= 12'h6af;
      20'h00466: out <= 12'h16d;
      20'h00467: out <= 12'h16d;
      20'h00468: out <= 12'h16d;
      20'h00469: out <= 12'h6af;
      20'h0046a: out <= 12'hfff;
      20'h0046b: out <= 12'h16d;
      20'h0046c: out <= 12'h222;
      20'h0046d: out <= 12'h222;
      20'h0046e: out <= 12'h222;
      20'h0046f: out <= 12'h222;
      20'h00470: out <= 12'h000;
      20'h00471: out <= 12'h000;
      20'h00472: out <= 12'h16d;
      20'h00473: out <= 12'hfff;
      20'h00474: out <= 12'h6af;
      20'h00475: out <= 12'h6af;
      20'h00476: out <= 12'h16d;
      20'h00477: out <= 12'h16d;
      20'h00478: out <= 12'h16d;
      20'h00479: out <= 12'h6af;
      20'h0047a: out <= 12'hfff;
      20'h0047b: out <= 12'h16d;
      20'h0047c: out <= 12'h000;
      20'h0047d: out <= 12'h000;
      20'h0047e: out <= 12'h000;
      20'h0047f: out <= 12'h000;
      20'h00480: out <= 12'h222;
      20'h00481: out <= 12'h6af;
      20'h00482: out <= 12'hfff;
      20'h00483: out <= 12'h6af;
      20'h00484: out <= 12'h222;
      20'h00485: out <= 12'h16d;
      20'h00486: out <= 12'h16d;
      20'h00487: out <= 12'h16d;
      20'h00488: out <= 12'hfff;
      20'h00489: out <= 12'h16d;
      20'h0048a: out <= 12'h16d;
      20'h0048b: out <= 12'h16d;
      20'h0048c: out <= 12'h222;
      20'h0048d: out <= 12'h6af;
      20'h0048e: out <= 12'hfff;
      20'h0048f: out <= 12'h6af;
      20'h00490: out <= 12'h000;
      20'h00491: out <= 12'h6af;
      20'h00492: out <= 12'h16d;
      20'h00493: out <= 12'h6af;
      20'h00494: out <= 12'h000;
      20'h00495: out <= 12'h16d;
      20'h00496: out <= 12'h16d;
      20'h00497: out <= 12'h16d;
      20'h00498: out <= 12'hfff;
      20'h00499: out <= 12'h16d;
      20'h0049a: out <= 12'h16d;
      20'h0049b: out <= 12'h16d;
      20'h0049c: out <= 12'h000;
      20'h0049d: out <= 12'h6af;
      20'h0049e: out <= 12'h16d;
      20'h0049f: out <= 12'h6af;
      20'h004a0: out <= 12'h222;
      20'h004a1: out <= 12'h222;
      20'h004a2: out <= 12'h222;
      20'h004a3: out <= 12'h222;
      20'h004a4: out <= 12'h16d;
      20'h004a5: out <= 12'hfff;
      20'h004a6: out <= 12'h6af;
      20'h004a7: out <= 12'h16d;
      20'h004a8: out <= 12'h16d;
      20'h004a9: out <= 12'h16d;
      20'h004aa: out <= 12'h6af;
      20'h004ab: out <= 12'h6af;
      20'h004ac: out <= 12'hfff;
      20'h004ad: out <= 12'h16d;
      20'h004ae: out <= 12'h222;
      20'h004af: out <= 12'h222;
      20'h004b0: out <= 12'h000;
      20'h004b1: out <= 12'h000;
      20'h004b2: out <= 12'h000;
      20'h004b3: out <= 12'h000;
      20'h004b4: out <= 12'h16d;
      20'h004b5: out <= 12'hfff;
      20'h004b6: out <= 12'h6af;
      20'h004b7: out <= 12'h16d;
      20'h004b8: out <= 12'h16d;
      20'h004b9: out <= 12'h16d;
      20'h004ba: out <= 12'h6af;
      20'h004bb: out <= 12'h6af;
      20'h004bc: out <= 12'hfff;
      20'h004bd: out <= 12'h16d;
      20'h004be: out <= 12'h000;
      20'h004bf: out <= 12'h000;
      20'h004c0: out <= 12'h222;
      20'h004c1: out <= 12'h6af;
      20'h004c2: out <= 12'h16d;
      20'h004c3: out <= 12'h16d;
      20'h004c4: out <= 12'hfff;
      20'h004c5: out <= 12'h6af;
      20'h004c6: out <= 12'h6af;
      20'h004c7: out <= 12'h16d;
      20'h004c8: out <= 12'h16d;
      20'h004c9: out <= 12'h16d;
      20'h004ca: out <= 12'h6af;
      20'h004cb: out <= 12'h6af;
      20'h004cc: out <= 12'hfff;
      20'h004cd: out <= 12'h16d;
      20'h004ce: out <= 12'h16d;
      20'h004cf: out <= 12'h6af;
      20'h004d0: out <= 12'h000;
      20'h004d1: out <= 12'h6af;
      20'h004d2: out <= 12'hfff;
      20'h004d3: out <= 12'h16d;
      20'h004d4: out <= 12'hfff;
      20'h004d5: out <= 12'h6af;
      20'h004d6: out <= 12'h6af;
      20'h004d7: out <= 12'h16d;
      20'h004d8: out <= 12'h16d;
      20'h004d9: out <= 12'h16d;
      20'h004da: out <= 12'h6af;
      20'h004db: out <= 12'h6af;
      20'h004dc: out <= 12'hfff;
      20'h004dd: out <= 12'h16d;
      20'h004de: out <= 12'hfff;
      20'h004df: out <= 12'h6af;
      20'h004e0: out <= 12'h603;
      20'h004e1: out <= 12'h603;
      20'h004e2: out <= 12'h603;
      20'h004e3: out <= 12'h603;
      20'h004e4: out <= 12'hb27;
      20'h004e5: out <= 12'hee9;
      20'h004e6: out <= 12'hee9;
      20'h004e7: out <= 12'hee9;
      20'h004e8: out <= 12'hee9;
      20'h004e9: out <= 12'hee9;
      20'h004ea: out <= 12'hee9;
      20'h004eb: out <= 12'hee9;
      20'h004ec: out <= 12'hb27;
      20'h004ed: out <= 12'hee9;
      20'h004ee: out <= 12'hee9;
      20'h004ef: out <= 12'hee9;
      20'h004f0: out <= 12'hee9;
      20'h004f1: out <= 12'hee9;
      20'h004f2: out <= 12'hee9;
      20'h004f3: out <= 12'hee9;
      20'h004f4: out <= 12'h000;
      20'h004f5: out <= 12'h000;
      20'h004f6: out <= 12'h000;
      20'h004f7: out <= 12'h000;
      20'h004f8: out <= 12'h000;
      20'h004f9: out <= 12'h000;
      20'h004fa: out <= 12'h000;
      20'h004fb: out <= 12'h000;
      20'h004fc: out <= 12'hb27;
      20'h004fd: out <= 12'hee9;
      20'h004fe: out <= 12'hee9;
      20'h004ff: out <= 12'hee9;
      20'h00500: out <= 12'hee9;
      20'h00501: out <= 12'hee9;
      20'h00502: out <= 12'hee9;
      20'h00503: out <= 12'hee9;
      20'h00504: out <= 12'h000;
      20'h00505: out <= 12'h000;
      20'h00506: out <= 12'h000;
      20'h00507: out <= 12'h000;
      20'h00508: out <= 12'h000;
      20'h00509: out <= 12'h000;
      20'h0050a: out <= 12'h000;
      20'h0050b: out <= 12'h000;
      20'h0050c: out <= 12'h000;
      20'h0050d: out <= 12'h000;
      20'h0050e: out <= 12'h000;
      20'h0050f: out <= 12'h000;
      20'h00510: out <= 12'h000;
      20'h00511: out <= 12'h000;
      20'h00512: out <= 12'h000;
      20'h00513: out <= 12'h000;
      20'h00514: out <= 12'hb27;
      20'h00515: out <= 12'hee9;
      20'h00516: out <= 12'hee9;
      20'h00517: out <= 12'hee9;
      20'h00518: out <= 12'hee9;
      20'h00519: out <= 12'hee9;
      20'h0051a: out <= 12'hee9;
      20'h0051b: out <= 12'hee9;
      20'h0051c: out <= 12'h000;
      20'h0051d: out <= 12'h000;
      20'h0051e: out <= 12'h000;
      20'h0051f: out <= 12'h000;
      20'h00520: out <= 12'h000;
      20'h00521: out <= 12'h000;
      20'h00522: out <= 12'h000;
      20'h00523: out <= 12'h000;
      20'h00524: out <= 12'hb27;
      20'h00525: out <= 12'hee9;
      20'h00526: out <= 12'hee9;
      20'h00527: out <= 12'hee9;
      20'h00528: out <= 12'hee9;
      20'h00529: out <= 12'hee9;
      20'h0052a: out <= 12'hee9;
      20'h0052b: out <= 12'hee9;
      20'h0052c: out <= 12'hb27;
      20'h0052d: out <= 12'hee9;
      20'h0052e: out <= 12'hee9;
      20'h0052f: out <= 12'hee9;
      20'h00530: out <= 12'hee9;
      20'h00531: out <= 12'hee9;
      20'h00532: out <= 12'hee9;
      20'h00533: out <= 12'hee9;
      20'h00534: out <= 12'h603;
      20'h00535: out <= 12'h603;
      20'h00536: out <= 12'h603;
      20'h00537: out <= 12'h603;
      20'h00538: out <= 12'hee9;
      20'h00539: out <= 12'hf87;
      20'h0053a: out <= 12'hee9;
      20'h0053b: out <= 12'hf87;
      20'h0053c: out <= 12'hf87;
      20'h0053d: out <= 12'hb27;
      20'h0053e: out <= 12'hf87;
      20'h0053f: out <= 12'hb27;
      20'h00540: out <= 12'hee9;
      20'h00541: out <= 12'hf87;
      20'h00542: out <= 12'hee9;
      20'h00543: out <= 12'hf87;
      20'h00544: out <= 12'hf87;
      20'h00545: out <= 12'hb27;
      20'h00546: out <= 12'hf87;
      20'h00547: out <= 12'hb27;
      20'h00548: out <= 12'hee9;
      20'h00549: out <= 12'hf87;
      20'h0054a: out <= 12'hee9;
      20'h0054b: out <= 12'hf87;
      20'h0054c: out <= 12'hf87;
      20'h0054d: out <= 12'hb27;
      20'h0054e: out <= 12'hf87;
      20'h0054f: out <= 12'hb27;
      20'h00550: out <= 12'hee9;
      20'h00551: out <= 12'hf87;
      20'h00552: out <= 12'hee9;
      20'h00553: out <= 12'hf87;
      20'h00554: out <= 12'hf87;
      20'h00555: out <= 12'hb27;
      20'h00556: out <= 12'hf87;
      20'h00557: out <= 12'hb27;
      20'h00558: out <= 12'hee9;
      20'h00559: out <= 12'hf87;
      20'h0055a: out <= 12'hee9;
      20'h0055b: out <= 12'hf87;
      20'h0055c: out <= 12'hf87;
      20'h0055d: out <= 12'hb27;
      20'h0055e: out <= 12'hf87;
      20'h0055f: out <= 12'hb27;
      20'h00560: out <= 12'hee9;
      20'h00561: out <= 12'hf87;
      20'h00562: out <= 12'hee9;
      20'h00563: out <= 12'hf87;
      20'h00564: out <= 12'hf87;
      20'h00565: out <= 12'hb27;
      20'h00566: out <= 12'hf87;
      20'h00567: out <= 12'hb27;
      20'h00568: out <= 12'hee9;
      20'h00569: out <= 12'hf87;
      20'h0056a: out <= 12'hee9;
      20'h0056b: out <= 12'hf87;
      20'h0056c: out <= 12'hf87;
      20'h0056d: out <= 12'hb27;
      20'h0056e: out <= 12'hf87;
      20'h0056f: out <= 12'hb27;
      20'h00570: out <= 12'hee9;
      20'h00571: out <= 12'hf87;
      20'h00572: out <= 12'hee9;
      20'h00573: out <= 12'hf87;
      20'h00574: out <= 12'hf87;
      20'h00575: out <= 12'hb27;
      20'h00576: out <= 12'hf87;
      20'h00577: out <= 12'hb27;
      20'h00578: out <= 12'h222;
      20'h00579: out <= 12'h222;
      20'h0057a: out <= 12'h16d;
      20'h0057b: out <= 12'h6af;
      20'h0057c: out <= 12'h6af;
      20'h0057d: out <= 12'h16d;
      20'h0057e: out <= 12'h16d;
      20'h0057f: out <= 12'h6af;
      20'h00580: out <= 12'h16d;
      20'h00581: out <= 12'h16d;
      20'h00582: out <= 12'h6af;
      20'h00583: out <= 12'h16d;
      20'h00584: out <= 12'h222;
      20'h00585: out <= 12'h222;
      20'h00586: out <= 12'h222;
      20'h00587: out <= 12'h222;
      20'h00588: out <= 12'h000;
      20'h00589: out <= 12'h000;
      20'h0058a: out <= 12'h16d;
      20'h0058b: out <= 12'h6af;
      20'h0058c: out <= 12'h6af;
      20'h0058d: out <= 12'h16d;
      20'h0058e: out <= 12'h16d;
      20'h0058f: out <= 12'h6af;
      20'h00590: out <= 12'h16d;
      20'h00591: out <= 12'h16d;
      20'h00592: out <= 12'h6af;
      20'h00593: out <= 12'h16d;
      20'h00594: out <= 12'h000;
      20'h00595: out <= 12'h000;
      20'h00596: out <= 12'h000;
      20'h00597: out <= 12'h000;
      20'h00598: out <= 12'h222;
      20'h00599: out <= 12'h6af;
      20'h0059a: out <= 12'h16d;
      20'h0059b: out <= 12'h16d;
      20'h0059c: out <= 12'h16d;
      20'h0059d: out <= 12'hfff;
      20'h0059e: out <= 12'h6af;
      20'h0059f: out <= 12'h16d;
      20'h005a0: out <= 12'h16d;
      20'h005a1: out <= 12'h16d;
      20'h005a2: out <= 12'h6af;
      20'h005a3: out <= 12'hfff;
      20'h005a4: out <= 12'h16d;
      20'h005a5: out <= 12'h16d;
      20'h005a6: out <= 12'h16d;
      20'h005a7: out <= 12'h6af;
      20'h005a8: out <= 12'h000;
      20'h005a9: out <= 12'h6af;
      20'h005aa: out <= 12'hfff;
      20'h005ab: out <= 12'h16d;
      20'h005ac: out <= 12'h16d;
      20'h005ad: out <= 12'hfff;
      20'h005ae: out <= 12'h6af;
      20'h005af: out <= 12'h16d;
      20'h005b0: out <= 12'h16d;
      20'h005b1: out <= 12'h16d;
      20'h005b2: out <= 12'h6af;
      20'h005b3: out <= 12'hfff;
      20'h005b4: out <= 12'h16d;
      20'h005b5: out <= 12'h16d;
      20'h005b6: out <= 12'hfff;
      20'h005b7: out <= 12'h6af;
      20'h005b8: out <= 12'h222;
      20'h005b9: out <= 12'h222;
      20'h005ba: out <= 12'h222;
      20'h005bb: out <= 12'h222;
      20'h005bc: out <= 12'h16d;
      20'h005bd: out <= 12'h6af;
      20'h005be: out <= 12'h16d;
      20'h005bf: out <= 12'h16d;
      20'h005c0: out <= 12'h6af;
      20'h005c1: out <= 12'h16d;
      20'h005c2: out <= 12'h16d;
      20'h005c3: out <= 12'h6af;
      20'h005c4: out <= 12'h6af;
      20'h005c5: out <= 12'h16d;
      20'h005c6: out <= 12'h222;
      20'h005c7: out <= 12'h222;
      20'h005c8: out <= 12'h000;
      20'h005c9: out <= 12'h000;
      20'h005ca: out <= 12'h000;
      20'h005cb: out <= 12'h000;
      20'h005cc: out <= 12'h16d;
      20'h005cd: out <= 12'h6af;
      20'h005ce: out <= 12'h16d;
      20'h005cf: out <= 12'h16d;
      20'h005d0: out <= 12'h6af;
      20'h005d1: out <= 12'h16d;
      20'h005d2: out <= 12'h16d;
      20'h005d3: out <= 12'h6af;
      20'h005d4: out <= 12'h6af;
      20'h005d5: out <= 12'h16d;
      20'h005d6: out <= 12'h000;
      20'h005d7: out <= 12'h000;
      20'h005d8: out <= 12'h222;
      20'h005d9: out <= 12'h6af;
      20'h005da: out <= 12'hfff;
      20'h005db: out <= 12'h16d;
      20'h005dc: out <= 12'h6af;
      20'h005dd: out <= 12'h6af;
      20'h005de: out <= 12'h16d;
      20'h005df: out <= 12'h16d;
      20'h005e0: out <= 12'h6af;
      20'h005e1: out <= 12'h16d;
      20'h005e2: out <= 12'h16d;
      20'h005e3: out <= 12'h6af;
      20'h005e4: out <= 12'h6af;
      20'h005e5: out <= 12'h16d;
      20'h005e6: out <= 12'hfff;
      20'h005e7: out <= 12'h6af;
      20'h005e8: out <= 12'h000;
      20'h005e9: out <= 12'h6af;
      20'h005ea: out <= 12'h16d;
      20'h005eb: out <= 12'h16d;
      20'h005ec: out <= 12'h6af;
      20'h005ed: out <= 12'h6af;
      20'h005ee: out <= 12'h16d;
      20'h005ef: out <= 12'h16d;
      20'h005f0: out <= 12'h6af;
      20'h005f1: out <= 12'h16d;
      20'h005f2: out <= 12'h16d;
      20'h005f3: out <= 12'h6af;
      20'h005f4: out <= 12'h6af;
      20'h005f5: out <= 12'h16d;
      20'h005f6: out <= 12'h16d;
      20'h005f7: out <= 12'h6af;
      20'h005f8: out <= 12'h603;
      20'h005f9: out <= 12'h603;
      20'h005fa: out <= 12'h603;
      20'h005fb: out <= 12'h603;
      20'h005fc: out <= 12'hb27;
      20'h005fd: out <= 12'hf87;
      20'h005fe: out <= 12'hf87;
      20'h005ff: out <= 12'hf87;
      20'h00600: out <= 12'hf87;
      20'h00601: out <= 12'hf87;
      20'h00602: out <= 12'hf87;
      20'h00603: out <= 12'hee9;
      20'h00604: out <= 12'hb27;
      20'h00605: out <= 12'hf87;
      20'h00606: out <= 12'hf87;
      20'h00607: out <= 12'hf87;
      20'h00608: out <= 12'hf87;
      20'h00609: out <= 12'hf87;
      20'h0060a: out <= 12'hf87;
      20'h0060b: out <= 12'hee9;
      20'h0060c: out <= 12'h000;
      20'h0060d: out <= 12'h000;
      20'h0060e: out <= 12'h000;
      20'h0060f: out <= 12'h000;
      20'h00610: out <= 12'h000;
      20'h00611: out <= 12'h000;
      20'h00612: out <= 12'h000;
      20'h00613: out <= 12'h000;
      20'h00614: out <= 12'hb27;
      20'h00615: out <= 12'hf87;
      20'h00616: out <= 12'hf87;
      20'h00617: out <= 12'hf87;
      20'h00618: out <= 12'hf87;
      20'h00619: out <= 12'hf87;
      20'h0061a: out <= 12'hf87;
      20'h0061b: out <= 12'hee9;
      20'h0061c: out <= 12'h000;
      20'h0061d: out <= 12'h000;
      20'h0061e: out <= 12'h000;
      20'h0061f: out <= 12'h000;
      20'h00620: out <= 12'h000;
      20'h00621: out <= 12'h000;
      20'h00622: out <= 12'h000;
      20'h00623: out <= 12'h000;
      20'h00624: out <= 12'h000;
      20'h00625: out <= 12'h000;
      20'h00626: out <= 12'h000;
      20'h00627: out <= 12'h000;
      20'h00628: out <= 12'h000;
      20'h00629: out <= 12'h000;
      20'h0062a: out <= 12'h000;
      20'h0062b: out <= 12'h000;
      20'h0062c: out <= 12'hb27;
      20'h0062d: out <= 12'hf87;
      20'h0062e: out <= 12'hf87;
      20'h0062f: out <= 12'hf87;
      20'h00630: out <= 12'hf87;
      20'h00631: out <= 12'hf87;
      20'h00632: out <= 12'hf87;
      20'h00633: out <= 12'hee9;
      20'h00634: out <= 12'h000;
      20'h00635: out <= 12'h000;
      20'h00636: out <= 12'h000;
      20'h00637: out <= 12'h000;
      20'h00638: out <= 12'h000;
      20'h00639: out <= 12'h000;
      20'h0063a: out <= 12'h000;
      20'h0063b: out <= 12'h000;
      20'h0063c: out <= 12'hb27;
      20'h0063d: out <= 12'hf87;
      20'h0063e: out <= 12'hf87;
      20'h0063f: out <= 12'hf87;
      20'h00640: out <= 12'hf87;
      20'h00641: out <= 12'hf87;
      20'h00642: out <= 12'hf87;
      20'h00643: out <= 12'hee9;
      20'h00644: out <= 12'hb27;
      20'h00645: out <= 12'hf87;
      20'h00646: out <= 12'hf87;
      20'h00647: out <= 12'hf87;
      20'h00648: out <= 12'hf87;
      20'h00649: out <= 12'hf87;
      20'h0064a: out <= 12'hf87;
      20'h0064b: out <= 12'hee9;
      20'h0064c: out <= 12'h603;
      20'h0064d: out <= 12'h603;
      20'h0064e: out <= 12'h603;
      20'h0064f: out <= 12'h603;
      20'h00650: out <= 12'hee9;
      20'h00651: out <= 12'hf87;
      20'h00652: out <= 12'hee9;
      20'h00653: out <= 12'hb27;
      20'h00654: out <= 12'hb27;
      20'h00655: out <= 12'hb27;
      20'h00656: out <= 12'hf87;
      20'h00657: out <= 12'hb27;
      20'h00658: out <= 12'hee9;
      20'h00659: out <= 12'hf87;
      20'h0065a: out <= 12'hee9;
      20'h0065b: out <= 12'hb27;
      20'h0065c: out <= 12'hb27;
      20'h0065d: out <= 12'hb27;
      20'h0065e: out <= 12'hf87;
      20'h0065f: out <= 12'hb27;
      20'h00660: out <= 12'hee9;
      20'h00661: out <= 12'hf87;
      20'h00662: out <= 12'hee9;
      20'h00663: out <= 12'hb27;
      20'h00664: out <= 12'hb27;
      20'h00665: out <= 12'hb27;
      20'h00666: out <= 12'hf87;
      20'h00667: out <= 12'hb27;
      20'h00668: out <= 12'hee9;
      20'h00669: out <= 12'hf87;
      20'h0066a: out <= 12'hee9;
      20'h0066b: out <= 12'hb27;
      20'h0066c: out <= 12'hb27;
      20'h0066d: out <= 12'hb27;
      20'h0066e: out <= 12'hf87;
      20'h0066f: out <= 12'hb27;
      20'h00670: out <= 12'hee9;
      20'h00671: out <= 12'hf87;
      20'h00672: out <= 12'hee9;
      20'h00673: out <= 12'hb27;
      20'h00674: out <= 12'hb27;
      20'h00675: out <= 12'hb27;
      20'h00676: out <= 12'hf87;
      20'h00677: out <= 12'hb27;
      20'h00678: out <= 12'hee9;
      20'h00679: out <= 12'hf87;
      20'h0067a: out <= 12'hee9;
      20'h0067b: out <= 12'hb27;
      20'h0067c: out <= 12'hb27;
      20'h0067d: out <= 12'hb27;
      20'h0067e: out <= 12'hf87;
      20'h0067f: out <= 12'hb27;
      20'h00680: out <= 12'hee9;
      20'h00681: out <= 12'hf87;
      20'h00682: out <= 12'hee9;
      20'h00683: out <= 12'hb27;
      20'h00684: out <= 12'hb27;
      20'h00685: out <= 12'hb27;
      20'h00686: out <= 12'hf87;
      20'h00687: out <= 12'hb27;
      20'h00688: out <= 12'hee9;
      20'h00689: out <= 12'hf87;
      20'h0068a: out <= 12'hee9;
      20'h0068b: out <= 12'hb27;
      20'h0068c: out <= 12'hb27;
      20'h0068d: out <= 12'hb27;
      20'h0068e: out <= 12'hf87;
      20'h0068f: out <= 12'hb27;
      20'h00690: out <= 12'h222;
      20'h00691: out <= 12'h222;
      20'h00692: out <= 12'h16d;
      20'h00693: out <= 12'h6af;
      20'h00694: out <= 12'h16d;
      20'h00695: out <= 12'h16d;
      20'h00696: out <= 12'h6af;
      20'h00697: out <= 12'hfff;
      20'h00698: out <= 12'h6af;
      20'h00699: out <= 12'h16d;
      20'h0069a: out <= 12'h16d;
      20'h0069b: out <= 12'h16d;
      20'h0069c: out <= 12'h16d;
      20'h0069d: out <= 12'h16d;
      20'h0069e: out <= 12'h16d;
      20'h0069f: out <= 12'h6af;
      20'h006a0: out <= 12'h000;
      20'h006a1: out <= 12'h000;
      20'h006a2: out <= 12'h16d;
      20'h006a3: out <= 12'h6af;
      20'h006a4: out <= 12'h16d;
      20'h006a5: out <= 12'h16d;
      20'h006a6: out <= 12'h6af;
      20'h006a7: out <= 12'hfff;
      20'h006a8: out <= 12'h6af;
      20'h006a9: out <= 12'h16d;
      20'h006aa: out <= 12'h16d;
      20'h006ab: out <= 12'h16d;
      20'h006ac: out <= 12'h16d;
      20'h006ad: out <= 12'h16d;
      20'h006ae: out <= 12'h16d;
      20'h006af: out <= 12'h6af;
      20'h006b0: out <= 12'h222;
      20'h006b1: out <= 12'h6af;
      20'h006b2: out <= 12'hfff;
      20'h006b3: out <= 12'h16d;
      20'h006b4: out <= 12'hfff;
      20'h006b5: out <= 12'h6af;
      20'h006b6: out <= 12'h16d;
      20'h006b7: out <= 12'h16d;
      20'h006b8: out <= 12'h6af;
      20'h006b9: out <= 12'h16d;
      20'h006ba: out <= 12'h16d;
      20'h006bb: out <= 12'h6af;
      20'h006bc: out <= 12'hfff;
      20'h006bd: out <= 12'h16d;
      20'h006be: out <= 12'hfff;
      20'h006bf: out <= 12'h6af;
      20'h006c0: out <= 12'h000;
      20'h006c1: out <= 12'h6af;
      20'h006c2: out <= 12'h16d;
      20'h006c3: out <= 12'h16d;
      20'h006c4: out <= 12'hfff;
      20'h006c5: out <= 12'h6af;
      20'h006c6: out <= 12'h16d;
      20'h006c7: out <= 12'h16d;
      20'h006c8: out <= 12'h6af;
      20'h006c9: out <= 12'h16d;
      20'h006ca: out <= 12'h16d;
      20'h006cb: out <= 12'h6af;
      20'h006cc: out <= 12'hfff;
      20'h006cd: out <= 12'h16d;
      20'h006ce: out <= 12'h16d;
      20'h006cf: out <= 12'h6af;
      20'h006d0: out <= 12'h6af;
      20'h006d1: out <= 12'h16d;
      20'h006d2: out <= 12'h16d;
      20'h006d3: out <= 12'h16d;
      20'h006d4: out <= 12'h16d;
      20'h006d5: out <= 12'h16d;
      20'h006d6: out <= 12'h16d;
      20'h006d7: out <= 12'h6af;
      20'h006d8: out <= 12'hfff;
      20'h006d9: out <= 12'h6af;
      20'h006da: out <= 12'h16d;
      20'h006db: out <= 12'h16d;
      20'h006dc: out <= 12'h6af;
      20'h006dd: out <= 12'h16d;
      20'h006de: out <= 12'h222;
      20'h006df: out <= 12'h222;
      20'h006e0: out <= 12'h6af;
      20'h006e1: out <= 12'h16d;
      20'h006e2: out <= 12'h16d;
      20'h006e3: out <= 12'h16d;
      20'h006e4: out <= 12'h16d;
      20'h006e5: out <= 12'h16d;
      20'h006e6: out <= 12'h16d;
      20'h006e7: out <= 12'h6af;
      20'h006e8: out <= 12'hfff;
      20'h006e9: out <= 12'h6af;
      20'h006ea: out <= 12'h16d;
      20'h006eb: out <= 12'h16d;
      20'h006ec: out <= 12'h6af;
      20'h006ed: out <= 12'h16d;
      20'h006ee: out <= 12'h000;
      20'h006ef: out <= 12'h000;
      20'h006f0: out <= 12'h222;
      20'h006f1: out <= 12'h6af;
      20'h006f2: out <= 12'h16d;
      20'h006f3: out <= 12'h16d;
      20'h006f4: out <= 12'h6af;
      20'h006f5: out <= 12'h16d;
      20'h006f6: out <= 12'h16d;
      20'h006f7: out <= 12'h6af;
      20'h006f8: out <= 12'hfff;
      20'h006f9: out <= 12'h6af;
      20'h006fa: out <= 12'h16d;
      20'h006fb: out <= 12'h16d;
      20'h006fc: out <= 12'h6af;
      20'h006fd: out <= 12'h16d;
      20'h006fe: out <= 12'h16d;
      20'h006ff: out <= 12'h6af;
      20'h00700: out <= 12'h000;
      20'h00701: out <= 12'h6af;
      20'h00702: out <= 12'hfff;
      20'h00703: out <= 12'h16d;
      20'h00704: out <= 12'h6af;
      20'h00705: out <= 12'h16d;
      20'h00706: out <= 12'h16d;
      20'h00707: out <= 12'h6af;
      20'h00708: out <= 12'hfff;
      20'h00709: out <= 12'h6af;
      20'h0070a: out <= 12'h16d;
      20'h0070b: out <= 12'h16d;
      20'h0070c: out <= 12'h6af;
      20'h0070d: out <= 12'h16d;
      20'h0070e: out <= 12'hfff;
      20'h0070f: out <= 12'h6af;
      20'h00710: out <= 12'h603;
      20'h00711: out <= 12'h603;
      20'h00712: out <= 12'h603;
      20'h00713: out <= 12'h603;
      20'h00714: out <= 12'hb27;
      20'h00715: out <= 12'hf87;
      20'h00716: out <= 12'hf87;
      20'h00717: out <= 12'hf87;
      20'h00718: out <= 12'hf87;
      20'h00719: out <= 12'hf87;
      20'h0071a: out <= 12'hf87;
      20'h0071b: out <= 12'hee9;
      20'h0071c: out <= 12'hb27;
      20'h0071d: out <= 12'hf87;
      20'h0071e: out <= 12'hf87;
      20'h0071f: out <= 12'hf87;
      20'h00720: out <= 12'hf87;
      20'h00721: out <= 12'hf87;
      20'h00722: out <= 12'hf87;
      20'h00723: out <= 12'hee9;
      20'h00724: out <= 12'h000;
      20'h00725: out <= 12'h000;
      20'h00726: out <= 12'h000;
      20'h00727: out <= 12'h000;
      20'h00728: out <= 12'h000;
      20'h00729: out <= 12'h000;
      20'h0072a: out <= 12'h000;
      20'h0072b: out <= 12'h000;
      20'h0072c: out <= 12'hb27;
      20'h0072d: out <= 12'hf87;
      20'h0072e: out <= 12'hf87;
      20'h0072f: out <= 12'hf87;
      20'h00730: out <= 12'hf87;
      20'h00731: out <= 12'hf87;
      20'h00732: out <= 12'hf87;
      20'h00733: out <= 12'hee9;
      20'h00734: out <= 12'h000;
      20'h00735: out <= 12'h000;
      20'h00736: out <= 12'h000;
      20'h00737: out <= 12'h000;
      20'h00738: out <= 12'h000;
      20'h00739: out <= 12'h000;
      20'h0073a: out <= 12'h000;
      20'h0073b: out <= 12'h000;
      20'h0073c: out <= 12'h000;
      20'h0073d: out <= 12'h000;
      20'h0073e: out <= 12'h000;
      20'h0073f: out <= 12'h000;
      20'h00740: out <= 12'h000;
      20'h00741: out <= 12'h000;
      20'h00742: out <= 12'h000;
      20'h00743: out <= 12'h000;
      20'h00744: out <= 12'hb27;
      20'h00745: out <= 12'hf87;
      20'h00746: out <= 12'hf87;
      20'h00747: out <= 12'hf87;
      20'h00748: out <= 12'hf87;
      20'h00749: out <= 12'hf87;
      20'h0074a: out <= 12'hf87;
      20'h0074b: out <= 12'hee9;
      20'h0074c: out <= 12'h000;
      20'h0074d: out <= 12'h000;
      20'h0074e: out <= 12'h000;
      20'h0074f: out <= 12'h000;
      20'h00750: out <= 12'h000;
      20'h00751: out <= 12'h000;
      20'h00752: out <= 12'h000;
      20'h00753: out <= 12'h000;
      20'h00754: out <= 12'hb27;
      20'h00755: out <= 12'hf87;
      20'h00756: out <= 12'hf87;
      20'h00757: out <= 12'hf87;
      20'h00758: out <= 12'hf87;
      20'h00759: out <= 12'hf87;
      20'h0075a: out <= 12'hf87;
      20'h0075b: out <= 12'hee9;
      20'h0075c: out <= 12'hb27;
      20'h0075d: out <= 12'hf87;
      20'h0075e: out <= 12'hf87;
      20'h0075f: out <= 12'hf87;
      20'h00760: out <= 12'hf87;
      20'h00761: out <= 12'hf87;
      20'h00762: out <= 12'hf87;
      20'h00763: out <= 12'hee9;
      20'h00764: out <= 12'h603;
      20'h00765: out <= 12'h603;
      20'h00766: out <= 12'h603;
      20'h00767: out <= 12'h603;
      20'h00768: out <= 12'hee9;
      20'h00769: out <= 12'hf87;
      20'h0076a: out <= 12'hf87;
      20'h0076b: out <= 12'hf87;
      20'h0076c: out <= 12'hf87;
      20'h0076d: out <= 12'hf87;
      20'h0076e: out <= 12'hf87;
      20'h0076f: out <= 12'hb27;
      20'h00770: out <= 12'hee9;
      20'h00771: out <= 12'hf87;
      20'h00772: out <= 12'hf87;
      20'h00773: out <= 12'hf87;
      20'h00774: out <= 12'hf87;
      20'h00775: out <= 12'hf87;
      20'h00776: out <= 12'hf87;
      20'h00777: out <= 12'hb27;
      20'h00778: out <= 12'hee9;
      20'h00779: out <= 12'hf87;
      20'h0077a: out <= 12'hf87;
      20'h0077b: out <= 12'hf87;
      20'h0077c: out <= 12'hf87;
      20'h0077d: out <= 12'hf87;
      20'h0077e: out <= 12'hf87;
      20'h0077f: out <= 12'hb27;
      20'h00780: out <= 12'hee9;
      20'h00781: out <= 12'hf87;
      20'h00782: out <= 12'hf87;
      20'h00783: out <= 12'hf87;
      20'h00784: out <= 12'hf87;
      20'h00785: out <= 12'hf87;
      20'h00786: out <= 12'hf87;
      20'h00787: out <= 12'hb27;
      20'h00788: out <= 12'hee9;
      20'h00789: out <= 12'hf87;
      20'h0078a: out <= 12'hf87;
      20'h0078b: out <= 12'hf87;
      20'h0078c: out <= 12'hf87;
      20'h0078d: out <= 12'hf87;
      20'h0078e: out <= 12'hf87;
      20'h0078f: out <= 12'hb27;
      20'h00790: out <= 12'hee9;
      20'h00791: out <= 12'hf87;
      20'h00792: out <= 12'hf87;
      20'h00793: out <= 12'hf87;
      20'h00794: out <= 12'hf87;
      20'h00795: out <= 12'hf87;
      20'h00796: out <= 12'hf87;
      20'h00797: out <= 12'hb27;
      20'h00798: out <= 12'hee9;
      20'h00799: out <= 12'hf87;
      20'h0079a: out <= 12'hf87;
      20'h0079b: out <= 12'hf87;
      20'h0079c: out <= 12'hf87;
      20'h0079d: out <= 12'hf87;
      20'h0079e: out <= 12'hf87;
      20'h0079f: out <= 12'hb27;
      20'h007a0: out <= 12'hee9;
      20'h007a1: out <= 12'hf87;
      20'h007a2: out <= 12'hf87;
      20'h007a3: out <= 12'hf87;
      20'h007a4: out <= 12'hf87;
      20'h007a5: out <= 12'hf87;
      20'h007a6: out <= 12'hf87;
      20'h007a7: out <= 12'hb27;
      20'h007a8: out <= 12'h222;
      20'h007a9: out <= 12'h222;
      20'h007aa: out <= 12'h16d;
      20'h007ab: out <= 12'h6af;
      20'h007ac: out <= 12'h16d;
      20'h007ad: out <= 12'h6af;
      20'h007ae: out <= 12'hfff;
      20'h007af: out <= 12'hfff;
      20'h007b0: out <= 12'hfff;
      20'h007b1: out <= 12'h6af;
      20'h007b2: out <= 12'h16d;
      20'h007b3: out <= 12'hfff;
      20'h007b4: out <= 12'hfff;
      20'h007b5: out <= 12'hfff;
      20'h007b6: out <= 12'hfff;
      20'h007b7: out <= 12'hfff;
      20'h007b8: out <= 12'h000;
      20'h007b9: out <= 12'h000;
      20'h007ba: out <= 12'h16d;
      20'h007bb: out <= 12'h6af;
      20'h007bc: out <= 12'h16d;
      20'h007bd: out <= 12'h6af;
      20'h007be: out <= 12'hfff;
      20'h007bf: out <= 12'hfff;
      20'h007c0: out <= 12'hfff;
      20'h007c1: out <= 12'h6af;
      20'h007c2: out <= 12'h16d;
      20'h007c3: out <= 12'hfff;
      20'h007c4: out <= 12'hfff;
      20'h007c5: out <= 12'hfff;
      20'h007c6: out <= 12'hfff;
      20'h007c7: out <= 12'hfff;
      20'h007c8: out <= 12'h222;
      20'h007c9: out <= 12'h6af;
      20'h007ca: out <= 12'h16d;
      20'h007cb: out <= 12'h16d;
      20'h007cc: out <= 12'h6af;
      20'h007cd: out <= 12'h16d;
      20'h007ce: out <= 12'h16d;
      20'h007cf: out <= 12'h6af;
      20'h007d0: out <= 12'hfff;
      20'h007d1: out <= 12'h6af;
      20'h007d2: out <= 12'h16d;
      20'h007d3: out <= 12'h16d;
      20'h007d4: out <= 12'h6af;
      20'h007d5: out <= 12'h16d;
      20'h007d6: out <= 12'h16d;
      20'h007d7: out <= 12'h6af;
      20'h007d8: out <= 12'h000;
      20'h007d9: out <= 12'h6af;
      20'h007da: out <= 12'hfff;
      20'h007db: out <= 12'h16d;
      20'h007dc: out <= 12'h6af;
      20'h007dd: out <= 12'h16d;
      20'h007de: out <= 12'h16d;
      20'h007df: out <= 12'h6af;
      20'h007e0: out <= 12'hfff;
      20'h007e1: out <= 12'h6af;
      20'h007e2: out <= 12'h16d;
      20'h007e3: out <= 12'h16d;
      20'h007e4: out <= 12'h6af;
      20'h007e5: out <= 12'h16d;
      20'h007e6: out <= 12'hfff;
      20'h007e7: out <= 12'h6af;
      20'h007e8: out <= 12'hfff;
      20'h007e9: out <= 12'hfff;
      20'h007ea: out <= 12'hfff;
      20'h007eb: out <= 12'hfff;
      20'h007ec: out <= 12'hfff;
      20'h007ed: out <= 12'h16d;
      20'h007ee: out <= 12'h6af;
      20'h007ef: out <= 12'hfff;
      20'h007f0: out <= 12'hfff;
      20'h007f1: out <= 12'hfff;
      20'h007f2: out <= 12'h6af;
      20'h007f3: out <= 12'h16d;
      20'h007f4: out <= 12'h6af;
      20'h007f5: out <= 12'h16d;
      20'h007f6: out <= 12'h222;
      20'h007f7: out <= 12'h222;
      20'h007f8: out <= 12'hfff;
      20'h007f9: out <= 12'hfff;
      20'h007fa: out <= 12'hfff;
      20'h007fb: out <= 12'hfff;
      20'h007fc: out <= 12'hfff;
      20'h007fd: out <= 12'h16d;
      20'h007fe: out <= 12'h6af;
      20'h007ff: out <= 12'hfff;
      20'h00800: out <= 12'hfff;
      20'h00801: out <= 12'hfff;
      20'h00802: out <= 12'h6af;
      20'h00803: out <= 12'h16d;
      20'h00804: out <= 12'h6af;
      20'h00805: out <= 12'h16d;
      20'h00806: out <= 12'h000;
      20'h00807: out <= 12'h000;
      20'h00808: out <= 12'h222;
      20'h00809: out <= 12'h6af;
      20'h0080a: out <= 12'hfff;
      20'h0080b: out <= 12'h16d;
      20'h0080c: out <= 12'h6af;
      20'h0080d: out <= 12'h16d;
      20'h0080e: out <= 12'h6af;
      20'h0080f: out <= 12'hfff;
      20'h00810: out <= 12'hfff;
      20'h00811: out <= 12'hfff;
      20'h00812: out <= 12'h6af;
      20'h00813: out <= 12'h16d;
      20'h00814: out <= 12'h6af;
      20'h00815: out <= 12'h16d;
      20'h00816: out <= 12'hfff;
      20'h00817: out <= 12'h6af;
      20'h00818: out <= 12'h000;
      20'h00819: out <= 12'h6af;
      20'h0081a: out <= 12'h16d;
      20'h0081b: out <= 12'h16d;
      20'h0081c: out <= 12'h6af;
      20'h0081d: out <= 12'h16d;
      20'h0081e: out <= 12'h6af;
      20'h0081f: out <= 12'hfff;
      20'h00820: out <= 12'hfff;
      20'h00821: out <= 12'hfff;
      20'h00822: out <= 12'h6af;
      20'h00823: out <= 12'h16d;
      20'h00824: out <= 12'h6af;
      20'h00825: out <= 12'h16d;
      20'h00826: out <= 12'h16d;
      20'h00827: out <= 12'h6af;
      20'h00828: out <= 12'h603;
      20'h00829: out <= 12'h603;
      20'h0082a: out <= 12'h603;
      20'h0082b: out <= 12'h603;
      20'h0082c: out <= 12'hb27;
      20'h0082d: out <= 12'hb27;
      20'h0082e: out <= 12'hb27;
      20'h0082f: out <= 12'hb27;
      20'h00830: out <= 12'hb27;
      20'h00831: out <= 12'hb27;
      20'h00832: out <= 12'hb27;
      20'h00833: out <= 12'hb27;
      20'h00834: out <= 12'hb27;
      20'h00835: out <= 12'hb27;
      20'h00836: out <= 12'hb27;
      20'h00837: out <= 12'hb27;
      20'h00838: out <= 12'hb27;
      20'h00839: out <= 12'hb27;
      20'h0083a: out <= 12'hb27;
      20'h0083b: out <= 12'hb27;
      20'h0083c: out <= 12'h000;
      20'h0083d: out <= 12'h000;
      20'h0083e: out <= 12'h000;
      20'h0083f: out <= 12'h000;
      20'h00840: out <= 12'h000;
      20'h00841: out <= 12'h000;
      20'h00842: out <= 12'h000;
      20'h00843: out <= 12'h000;
      20'h00844: out <= 12'hb27;
      20'h00845: out <= 12'hb27;
      20'h00846: out <= 12'hb27;
      20'h00847: out <= 12'hb27;
      20'h00848: out <= 12'hb27;
      20'h00849: out <= 12'hb27;
      20'h0084a: out <= 12'hb27;
      20'h0084b: out <= 12'hb27;
      20'h0084c: out <= 12'h000;
      20'h0084d: out <= 12'h000;
      20'h0084e: out <= 12'h000;
      20'h0084f: out <= 12'h000;
      20'h00850: out <= 12'h000;
      20'h00851: out <= 12'h000;
      20'h00852: out <= 12'h000;
      20'h00853: out <= 12'h000;
      20'h00854: out <= 12'h000;
      20'h00855: out <= 12'h000;
      20'h00856: out <= 12'h000;
      20'h00857: out <= 12'h000;
      20'h00858: out <= 12'h000;
      20'h00859: out <= 12'h000;
      20'h0085a: out <= 12'h000;
      20'h0085b: out <= 12'h000;
      20'h0085c: out <= 12'hb27;
      20'h0085d: out <= 12'hb27;
      20'h0085e: out <= 12'hb27;
      20'h0085f: out <= 12'hb27;
      20'h00860: out <= 12'hb27;
      20'h00861: out <= 12'hb27;
      20'h00862: out <= 12'hb27;
      20'h00863: out <= 12'hb27;
      20'h00864: out <= 12'h000;
      20'h00865: out <= 12'h000;
      20'h00866: out <= 12'h000;
      20'h00867: out <= 12'h000;
      20'h00868: out <= 12'h000;
      20'h00869: out <= 12'h000;
      20'h0086a: out <= 12'h000;
      20'h0086b: out <= 12'h000;
      20'h0086c: out <= 12'hb27;
      20'h0086d: out <= 12'hb27;
      20'h0086e: out <= 12'hb27;
      20'h0086f: out <= 12'hb27;
      20'h00870: out <= 12'hb27;
      20'h00871: out <= 12'hb27;
      20'h00872: out <= 12'hb27;
      20'h00873: out <= 12'hb27;
      20'h00874: out <= 12'hb27;
      20'h00875: out <= 12'hb27;
      20'h00876: out <= 12'hb27;
      20'h00877: out <= 12'hb27;
      20'h00878: out <= 12'hb27;
      20'h00879: out <= 12'hb27;
      20'h0087a: out <= 12'hb27;
      20'h0087b: out <= 12'hb27;
      20'h0087c: out <= 12'h603;
      20'h0087d: out <= 12'h603;
      20'h0087e: out <= 12'h603;
      20'h0087f: out <= 12'h603;
      20'h00880: out <= 12'hb27;
      20'h00881: out <= 12'hb27;
      20'h00882: out <= 12'hb27;
      20'h00883: out <= 12'hb27;
      20'h00884: out <= 12'hb27;
      20'h00885: out <= 12'hb27;
      20'h00886: out <= 12'hb27;
      20'h00887: out <= 12'hb27;
      20'h00888: out <= 12'hb27;
      20'h00889: out <= 12'hb27;
      20'h0088a: out <= 12'hb27;
      20'h0088b: out <= 12'hb27;
      20'h0088c: out <= 12'hb27;
      20'h0088d: out <= 12'hb27;
      20'h0088e: out <= 12'hb27;
      20'h0088f: out <= 12'hb27;
      20'h00890: out <= 12'hb27;
      20'h00891: out <= 12'hb27;
      20'h00892: out <= 12'hb27;
      20'h00893: out <= 12'hb27;
      20'h00894: out <= 12'hb27;
      20'h00895: out <= 12'hb27;
      20'h00896: out <= 12'hb27;
      20'h00897: out <= 12'hb27;
      20'h00898: out <= 12'hb27;
      20'h00899: out <= 12'hb27;
      20'h0089a: out <= 12'hb27;
      20'h0089b: out <= 12'hb27;
      20'h0089c: out <= 12'hb27;
      20'h0089d: out <= 12'hb27;
      20'h0089e: out <= 12'hb27;
      20'h0089f: out <= 12'hb27;
      20'h008a0: out <= 12'hb27;
      20'h008a1: out <= 12'hb27;
      20'h008a2: out <= 12'hb27;
      20'h008a3: out <= 12'hb27;
      20'h008a4: out <= 12'hb27;
      20'h008a5: out <= 12'hb27;
      20'h008a6: out <= 12'hb27;
      20'h008a7: out <= 12'hb27;
      20'h008a8: out <= 12'hb27;
      20'h008a9: out <= 12'hb27;
      20'h008aa: out <= 12'hb27;
      20'h008ab: out <= 12'hb27;
      20'h008ac: out <= 12'hb27;
      20'h008ad: out <= 12'hb27;
      20'h008ae: out <= 12'hb27;
      20'h008af: out <= 12'hb27;
      20'h008b0: out <= 12'hb27;
      20'h008b1: out <= 12'hb27;
      20'h008b2: out <= 12'hb27;
      20'h008b3: out <= 12'hb27;
      20'h008b4: out <= 12'hb27;
      20'h008b5: out <= 12'hb27;
      20'h008b6: out <= 12'hb27;
      20'h008b7: out <= 12'hb27;
      20'h008b8: out <= 12'hb27;
      20'h008b9: out <= 12'hb27;
      20'h008ba: out <= 12'hb27;
      20'h008bb: out <= 12'hb27;
      20'h008bc: out <= 12'hb27;
      20'h008bd: out <= 12'hb27;
      20'h008be: out <= 12'hb27;
      20'h008bf: out <= 12'hb27;
      20'h008c0: out <= 12'h222;
      20'h008c1: out <= 12'h222;
      20'h008c2: out <= 12'h16d;
      20'h008c3: out <= 12'h6af;
      20'h008c4: out <= 12'h16d;
      20'h008c5: out <= 12'h16d;
      20'h008c6: out <= 12'h6af;
      20'h008c7: out <= 12'hfff;
      20'h008c8: out <= 12'h6af;
      20'h008c9: out <= 12'h16d;
      20'h008ca: out <= 12'h16d;
      20'h008cb: out <= 12'h16d;
      20'h008cc: out <= 12'h16d;
      20'h008cd: out <= 12'h16d;
      20'h008ce: out <= 12'h16d;
      20'h008cf: out <= 12'h6af;
      20'h008d0: out <= 12'h000;
      20'h008d1: out <= 12'h000;
      20'h008d2: out <= 12'h16d;
      20'h008d3: out <= 12'h6af;
      20'h008d4: out <= 12'h16d;
      20'h008d5: out <= 12'h16d;
      20'h008d6: out <= 12'h6af;
      20'h008d7: out <= 12'hfff;
      20'h008d8: out <= 12'h6af;
      20'h008d9: out <= 12'h16d;
      20'h008da: out <= 12'h16d;
      20'h008db: out <= 12'h16d;
      20'h008dc: out <= 12'h16d;
      20'h008dd: out <= 12'h16d;
      20'h008de: out <= 12'h16d;
      20'h008df: out <= 12'h6af;
      20'h008e0: out <= 12'h222;
      20'h008e1: out <= 12'h6af;
      20'h008e2: out <= 12'hfff;
      20'h008e3: out <= 12'h16d;
      20'h008e4: out <= 12'h6af;
      20'h008e5: out <= 12'h16d;
      20'h008e6: out <= 12'h6af;
      20'h008e7: out <= 12'hfff;
      20'h008e8: out <= 12'hfff;
      20'h008e9: out <= 12'hfff;
      20'h008ea: out <= 12'h6af;
      20'h008eb: out <= 12'h16d;
      20'h008ec: out <= 12'h6af;
      20'h008ed: out <= 12'h16d;
      20'h008ee: out <= 12'hfff;
      20'h008ef: out <= 12'h6af;
      20'h008f0: out <= 12'h000;
      20'h008f1: out <= 12'h6af;
      20'h008f2: out <= 12'h16d;
      20'h008f3: out <= 12'h16d;
      20'h008f4: out <= 12'h6af;
      20'h008f5: out <= 12'h16d;
      20'h008f6: out <= 12'h6af;
      20'h008f7: out <= 12'hfff;
      20'h008f8: out <= 12'hfff;
      20'h008f9: out <= 12'hfff;
      20'h008fa: out <= 12'h6af;
      20'h008fb: out <= 12'h16d;
      20'h008fc: out <= 12'h6af;
      20'h008fd: out <= 12'h16d;
      20'h008fe: out <= 12'h16d;
      20'h008ff: out <= 12'h6af;
      20'h00900: out <= 12'h6af;
      20'h00901: out <= 12'h16d;
      20'h00902: out <= 12'h16d;
      20'h00903: out <= 12'h16d;
      20'h00904: out <= 12'h16d;
      20'h00905: out <= 12'h16d;
      20'h00906: out <= 12'h16d;
      20'h00907: out <= 12'h6af;
      20'h00908: out <= 12'hfff;
      20'h00909: out <= 12'h6af;
      20'h0090a: out <= 12'h16d;
      20'h0090b: out <= 12'h16d;
      20'h0090c: out <= 12'h6af;
      20'h0090d: out <= 12'h16d;
      20'h0090e: out <= 12'h222;
      20'h0090f: out <= 12'h222;
      20'h00910: out <= 12'h6af;
      20'h00911: out <= 12'h16d;
      20'h00912: out <= 12'h16d;
      20'h00913: out <= 12'h16d;
      20'h00914: out <= 12'h16d;
      20'h00915: out <= 12'h16d;
      20'h00916: out <= 12'h16d;
      20'h00917: out <= 12'h6af;
      20'h00918: out <= 12'hfff;
      20'h00919: out <= 12'h6af;
      20'h0091a: out <= 12'h16d;
      20'h0091b: out <= 12'h16d;
      20'h0091c: out <= 12'h6af;
      20'h0091d: out <= 12'h16d;
      20'h0091e: out <= 12'h000;
      20'h0091f: out <= 12'h000;
      20'h00920: out <= 12'h222;
      20'h00921: out <= 12'h6af;
      20'h00922: out <= 12'h16d;
      20'h00923: out <= 12'h16d;
      20'h00924: out <= 12'h6af;
      20'h00925: out <= 12'h16d;
      20'h00926: out <= 12'h16d;
      20'h00927: out <= 12'h6af;
      20'h00928: out <= 12'hfff;
      20'h00929: out <= 12'h6af;
      20'h0092a: out <= 12'h16d;
      20'h0092b: out <= 12'h16d;
      20'h0092c: out <= 12'h6af;
      20'h0092d: out <= 12'h16d;
      20'h0092e: out <= 12'h16d;
      20'h0092f: out <= 12'h6af;
      20'h00930: out <= 12'h000;
      20'h00931: out <= 12'h6af;
      20'h00932: out <= 12'hfff;
      20'h00933: out <= 12'h16d;
      20'h00934: out <= 12'h6af;
      20'h00935: out <= 12'h16d;
      20'h00936: out <= 12'h16d;
      20'h00937: out <= 12'h6af;
      20'h00938: out <= 12'hfff;
      20'h00939: out <= 12'h6af;
      20'h0093a: out <= 12'h16d;
      20'h0093b: out <= 12'h16d;
      20'h0093c: out <= 12'h6af;
      20'h0093d: out <= 12'h16d;
      20'h0093e: out <= 12'hfff;
      20'h0093f: out <= 12'h6af;
      20'h00940: out <= 12'h603;
      20'h00941: out <= 12'h603;
      20'h00942: out <= 12'h603;
      20'h00943: out <= 12'h603;
      20'h00944: out <= 12'hee9;
      20'h00945: out <= 12'hee9;
      20'h00946: out <= 12'hee9;
      20'h00947: out <= 12'hee9;
      20'h00948: out <= 12'hb27;
      20'h00949: out <= 12'hee9;
      20'h0094a: out <= 12'hee9;
      20'h0094b: out <= 12'hee9;
      20'h0094c: out <= 12'hee9;
      20'h0094d: out <= 12'hee9;
      20'h0094e: out <= 12'hee9;
      20'h0094f: out <= 12'hee9;
      20'h00950: out <= 12'hb27;
      20'h00951: out <= 12'hee9;
      20'h00952: out <= 12'hee9;
      20'h00953: out <= 12'hee9;
      20'h00954: out <= 12'h000;
      20'h00955: out <= 12'h000;
      20'h00956: out <= 12'h000;
      20'h00957: out <= 12'h000;
      20'h00958: out <= 12'h000;
      20'h00959: out <= 12'h000;
      20'h0095a: out <= 12'h000;
      20'h0095b: out <= 12'h000;
      20'h0095c: out <= 12'hee9;
      20'h0095d: out <= 12'hee9;
      20'h0095e: out <= 12'hee9;
      20'h0095f: out <= 12'hee9;
      20'h00960: out <= 12'hb27;
      20'h00961: out <= 12'hee9;
      20'h00962: out <= 12'hee9;
      20'h00963: out <= 12'hee9;
      20'h00964: out <= 12'hee9;
      20'h00965: out <= 12'hee9;
      20'h00966: out <= 12'hee9;
      20'h00967: out <= 12'hee9;
      20'h00968: out <= 12'hb27;
      20'h00969: out <= 12'hee9;
      20'h0096a: out <= 12'hee9;
      20'h0096b: out <= 12'hee9;
      20'h0096c: out <= 12'hee9;
      20'h0096d: out <= 12'hee9;
      20'h0096e: out <= 12'hee9;
      20'h0096f: out <= 12'hee9;
      20'h00970: out <= 12'hb27;
      20'h00971: out <= 12'hee9;
      20'h00972: out <= 12'hee9;
      20'h00973: out <= 12'hee9;
      20'h00974: out <= 12'hee9;
      20'h00975: out <= 12'hee9;
      20'h00976: out <= 12'hee9;
      20'h00977: out <= 12'hee9;
      20'h00978: out <= 12'hb27;
      20'h00979: out <= 12'hee9;
      20'h0097a: out <= 12'hee9;
      20'h0097b: out <= 12'hee9;
      20'h0097c: out <= 12'h000;
      20'h0097d: out <= 12'h000;
      20'h0097e: out <= 12'h000;
      20'h0097f: out <= 12'h000;
      20'h00980: out <= 12'h000;
      20'h00981: out <= 12'h000;
      20'h00982: out <= 12'h000;
      20'h00983: out <= 12'h000;
      20'h00984: out <= 12'h000;
      20'h00985: out <= 12'h000;
      20'h00986: out <= 12'h000;
      20'h00987: out <= 12'h000;
      20'h00988: out <= 12'h000;
      20'h00989: out <= 12'h000;
      20'h0098a: out <= 12'h000;
      20'h0098b: out <= 12'h000;
      20'h0098c: out <= 12'h000;
      20'h0098d: out <= 12'h000;
      20'h0098e: out <= 12'h000;
      20'h0098f: out <= 12'h000;
      20'h00990: out <= 12'h000;
      20'h00991: out <= 12'h000;
      20'h00992: out <= 12'h000;
      20'h00993: out <= 12'h000;
      20'h00994: out <= 12'h603;
      20'h00995: out <= 12'h603;
      20'h00996: out <= 12'h603;
      20'h00997: out <= 12'h603;
      20'h00998: out <= 12'hee9;
      20'h00999: out <= 12'hee9;
      20'h0099a: out <= 12'hee9;
      20'h0099b: out <= 12'hee9;
      20'h0099c: out <= 12'hee9;
      20'h0099d: out <= 12'hee9;
      20'h0099e: out <= 12'hee9;
      20'h0099f: out <= 12'hb27;
      20'h009a0: out <= 12'h000;
      20'h009a1: out <= 12'h000;
      20'h009a2: out <= 12'h000;
      20'h009a3: out <= 12'h000;
      20'h009a4: out <= 12'h000;
      20'h009a5: out <= 12'h000;
      20'h009a6: out <= 12'h000;
      20'h009a7: out <= 12'h000;
      20'h009a8: out <= 12'h000;
      20'h009a9: out <= 12'h000;
      20'h009aa: out <= 12'h000;
      20'h009ab: out <= 12'h000;
      20'h009ac: out <= 12'h000;
      20'h009ad: out <= 12'h000;
      20'h009ae: out <= 12'h000;
      20'h009af: out <= 12'h000;
      20'h009b0: out <= 12'h000;
      20'h009b1: out <= 12'h000;
      20'h009b2: out <= 12'h000;
      20'h009b3: out <= 12'h000;
      20'h009b4: out <= 12'h000;
      20'h009b5: out <= 12'h000;
      20'h009b6: out <= 12'h000;
      20'h009b7: out <= 12'h000;
      20'h009b8: out <= 12'h000;
      20'h009b9: out <= 12'h000;
      20'h009ba: out <= 12'h000;
      20'h009bb: out <= 12'h000;
      20'h009bc: out <= 12'h000;
      20'h009bd: out <= 12'h000;
      20'h009be: out <= 12'h000;
      20'h009bf: out <= 12'h000;
      20'h009c0: out <= 12'h000;
      20'h009c1: out <= 12'h000;
      20'h009c2: out <= 12'h000;
      20'h009c3: out <= 12'h000;
      20'h009c4: out <= 12'h000;
      20'h009c5: out <= 12'h000;
      20'h009c6: out <= 12'h000;
      20'h009c7: out <= 12'h000;
      20'h009c8: out <= 12'h000;
      20'h009c9: out <= 12'h000;
      20'h009ca: out <= 12'h000;
      20'h009cb: out <= 12'h000;
      20'h009cc: out <= 12'h000;
      20'h009cd: out <= 12'h000;
      20'h009ce: out <= 12'h000;
      20'h009cf: out <= 12'h000;
      20'h009d0: out <= 12'h000;
      20'h009d1: out <= 12'h000;
      20'h009d2: out <= 12'h000;
      20'h009d3: out <= 12'h000;
      20'h009d4: out <= 12'h000;
      20'h009d5: out <= 12'h000;
      20'h009d6: out <= 12'h000;
      20'h009d7: out <= 12'h000;
      20'h009d8: out <= 12'h222;
      20'h009d9: out <= 12'h222;
      20'h009da: out <= 12'h16d;
      20'h009db: out <= 12'h6af;
      20'h009dc: out <= 12'h6af;
      20'h009dd: out <= 12'h16d;
      20'h009de: out <= 12'h16d;
      20'h009df: out <= 12'h6af;
      20'h009e0: out <= 12'h16d;
      20'h009e1: out <= 12'h16d;
      20'h009e2: out <= 12'h6af;
      20'h009e3: out <= 12'h16d;
      20'h009e4: out <= 12'h222;
      20'h009e5: out <= 12'h222;
      20'h009e6: out <= 12'h222;
      20'h009e7: out <= 12'h222;
      20'h009e8: out <= 12'h000;
      20'h009e9: out <= 12'h000;
      20'h009ea: out <= 12'h16d;
      20'h009eb: out <= 12'h6af;
      20'h009ec: out <= 12'h6af;
      20'h009ed: out <= 12'h16d;
      20'h009ee: out <= 12'h16d;
      20'h009ef: out <= 12'h6af;
      20'h009f0: out <= 12'h16d;
      20'h009f1: out <= 12'h16d;
      20'h009f2: out <= 12'h6af;
      20'h009f3: out <= 12'h16d;
      20'h009f4: out <= 12'h000;
      20'h009f5: out <= 12'h000;
      20'h009f6: out <= 12'h000;
      20'h009f7: out <= 12'h000;
      20'h009f8: out <= 12'h222;
      20'h009f9: out <= 12'h6af;
      20'h009fa: out <= 12'h16d;
      20'h009fb: out <= 12'h16d;
      20'h009fc: out <= 12'h6af;
      20'h009fd: out <= 12'h16d;
      20'h009fe: out <= 12'h16d;
      20'h009ff: out <= 12'h6af;
      20'h00a00: out <= 12'hfff;
      20'h00a01: out <= 12'h6af;
      20'h00a02: out <= 12'h16d;
      20'h00a03: out <= 12'h16d;
      20'h00a04: out <= 12'h6af;
      20'h00a05: out <= 12'h16d;
      20'h00a06: out <= 12'h16d;
      20'h00a07: out <= 12'h6af;
      20'h00a08: out <= 12'h000;
      20'h00a09: out <= 12'h6af;
      20'h00a0a: out <= 12'hfff;
      20'h00a0b: out <= 12'h16d;
      20'h00a0c: out <= 12'h6af;
      20'h00a0d: out <= 12'h16d;
      20'h00a0e: out <= 12'h16d;
      20'h00a0f: out <= 12'h6af;
      20'h00a10: out <= 12'hfff;
      20'h00a11: out <= 12'h6af;
      20'h00a12: out <= 12'h16d;
      20'h00a13: out <= 12'h16d;
      20'h00a14: out <= 12'h6af;
      20'h00a15: out <= 12'h16d;
      20'h00a16: out <= 12'hfff;
      20'h00a17: out <= 12'h6af;
      20'h00a18: out <= 12'h222;
      20'h00a19: out <= 12'h222;
      20'h00a1a: out <= 12'h222;
      20'h00a1b: out <= 12'h222;
      20'h00a1c: out <= 12'h16d;
      20'h00a1d: out <= 12'h6af;
      20'h00a1e: out <= 12'h16d;
      20'h00a1f: out <= 12'h16d;
      20'h00a20: out <= 12'h6af;
      20'h00a21: out <= 12'h16d;
      20'h00a22: out <= 12'h16d;
      20'h00a23: out <= 12'h6af;
      20'h00a24: out <= 12'h6af;
      20'h00a25: out <= 12'h16d;
      20'h00a26: out <= 12'h222;
      20'h00a27: out <= 12'h222;
      20'h00a28: out <= 12'h000;
      20'h00a29: out <= 12'h000;
      20'h00a2a: out <= 12'h000;
      20'h00a2b: out <= 12'h000;
      20'h00a2c: out <= 12'h16d;
      20'h00a2d: out <= 12'h6af;
      20'h00a2e: out <= 12'h16d;
      20'h00a2f: out <= 12'h16d;
      20'h00a30: out <= 12'h6af;
      20'h00a31: out <= 12'h16d;
      20'h00a32: out <= 12'h16d;
      20'h00a33: out <= 12'h6af;
      20'h00a34: out <= 12'h6af;
      20'h00a35: out <= 12'h16d;
      20'h00a36: out <= 12'h000;
      20'h00a37: out <= 12'h000;
      20'h00a38: out <= 12'h222;
      20'h00a39: out <= 12'h6af;
      20'h00a3a: out <= 12'hfff;
      20'h00a3b: out <= 12'h16d;
      20'h00a3c: out <= 12'hfff;
      20'h00a3d: out <= 12'h6af;
      20'h00a3e: out <= 12'h16d;
      20'h00a3f: out <= 12'h16d;
      20'h00a40: out <= 12'h6af;
      20'h00a41: out <= 12'h16d;
      20'h00a42: out <= 12'h16d;
      20'h00a43: out <= 12'h6af;
      20'h00a44: out <= 12'hfff;
      20'h00a45: out <= 12'h16d;
      20'h00a46: out <= 12'hfff;
      20'h00a47: out <= 12'h6af;
      20'h00a48: out <= 12'h000;
      20'h00a49: out <= 12'h6af;
      20'h00a4a: out <= 12'h16d;
      20'h00a4b: out <= 12'h16d;
      20'h00a4c: out <= 12'hfff;
      20'h00a4d: out <= 12'h6af;
      20'h00a4e: out <= 12'h16d;
      20'h00a4f: out <= 12'h16d;
      20'h00a50: out <= 12'h6af;
      20'h00a51: out <= 12'h16d;
      20'h00a52: out <= 12'h16d;
      20'h00a53: out <= 12'h6af;
      20'h00a54: out <= 12'hfff;
      20'h00a55: out <= 12'h16d;
      20'h00a56: out <= 12'h16d;
      20'h00a57: out <= 12'h6af;
      20'h00a58: out <= 12'h603;
      20'h00a59: out <= 12'h603;
      20'h00a5a: out <= 12'h603;
      20'h00a5b: out <= 12'h603;
      20'h00a5c: out <= 12'hf87;
      20'h00a5d: out <= 12'hf87;
      20'h00a5e: out <= 12'hf87;
      20'h00a5f: out <= 12'hee9;
      20'h00a60: out <= 12'hb27;
      20'h00a61: out <= 12'hf87;
      20'h00a62: out <= 12'hf87;
      20'h00a63: out <= 12'hf87;
      20'h00a64: out <= 12'hf87;
      20'h00a65: out <= 12'hf87;
      20'h00a66: out <= 12'hf87;
      20'h00a67: out <= 12'hee9;
      20'h00a68: out <= 12'hb27;
      20'h00a69: out <= 12'hf87;
      20'h00a6a: out <= 12'hf87;
      20'h00a6b: out <= 12'hf87;
      20'h00a6c: out <= 12'h000;
      20'h00a6d: out <= 12'h000;
      20'h00a6e: out <= 12'h000;
      20'h00a6f: out <= 12'h000;
      20'h00a70: out <= 12'h000;
      20'h00a71: out <= 12'h000;
      20'h00a72: out <= 12'h000;
      20'h00a73: out <= 12'h000;
      20'h00a74: out <= 12'hf87;
      20'h00a75: out <= 12'hf87;
      20'h00a76: out <= 12'hf87;
      20'h00a77: out <= 12'hee9;
      20'h00a78: out <= 12'hb27;
      20'h00a79: out <= 12'hf87;
      20'h00a7a: out <= 12'hf87;
      20'h00a7b: out <= 12'hf87;
      20'h00a7c: out <= 12'hf87;
      20'h00a7d: out <= 12'hf87;
      20'h00a7e: out <= 12'hf87;
      20'h00a7f: out <= 12'hee9;
      20'h00a80: out <= 12'hb27;
      20'h00a81: out <= 12'hf87;
      20'h00a82: out <= 12'hf87;
      20'h00a83: out <= 12'hf87;
      20'h00a84: out <= 12'hf87;
      20'h00a85: out <= 12'hf87;
      20'h00a86: out <= 12'hf87;
      20'h00a87: out <= 12'hee9;
      20'h00a88: out <= 12'hb27;
      20'h00a89: out <= 12'hf87;
      20'h00a8a: out <= 12'hf87;
      20'h00a8b: out <= 12'hf87;
      20'h00a8c: out <= 12'hf87;
      20'h00a8d: out <= 12'hf87;
      20'h00a8e: out <= 12'hf87;
      20'h00a8f: out <= 12'hee9;
      20'h00a90: out <= 12'hb27;
      20'h00a91: out <= 12'hf87;
      20'h00a92: out <= 12'hf87;
      20'h00a93: out <= 12'hf87;
      20'h00a94: out <= 12'h000;
      20'h00a95: out <= 12'h000;
      20'h00a96: out <= 12'h000;
      20'h00a97: out <= 12'h000;
      20'h00a98: out <= 12'h000;
      20'h00a99: out <= 12'h000;
      20'h00a9a: out <= 12'h000;
      20'h00a9b: out <= 12'h000;
      20'h00a9c: out <= 12'h000;
      20'h00a9d: out <= 12'h000;
      20'h00a9e: out <= 12'h000;
      20'h00a9f: out <= 12'h000;
      20'h00aa0: out <= 12'h000;
      20'h00aa1: out <= 12'h000;
      20'h00aa2: out <= 12'h000;
      20'h00aa3: out <= 12'h000;
      20'h00aa4: out <= 12'h000;
      20'h00aa5: out <= 12'h000;
      20'h00aa6: out <= 12'h000;
      20'h00aa7: out <= 12'h000;
      20'h00aa8: out <= 12'h000;
      20'h00aa9: out <= 12'h000;
      20'h00aaa: out <= 12'h000;
      20'h00aab: out <= 12'h000;
      20'h00aac: out <= 12'h603;
      20'h00aad: out <= 12'h603;
      20'h00aae: out <= 12'h603;
      20'h00aaf: out <= 12'h603;
      20'h00ab0: out <= 12'hee9;
      20'h00ab1: out <= 12'hf87;
      20'h00ab2: out <= 12'hf87;
      20'h00ab3: out <= 12'hf87;
      20'h00ab4: out <= 12'hf87;
      20'h00ab5: out <= 12'hf87;
      20'h00ab6: out <= 12'hf87;
      20'h00ab7: out <= 12'hb27;
      20'h00ab8: out <= 12'h000;
      20'h00ab9: out <= 12'h000;
      20'h00aba: out <= 12'h000;
      20'h00abb: out <= 12'h000;
      20'h00abc: out <= 12'h000;
      20'h00abd: out <= 12'h000;
      20'h00abe: out <= 12'h000;
      20'h00abf: out <= 12'h000;
      20'h00ac0: out <= 12'h000;
      20'h00ac1: out <= 12'h000;
      20'h00ac2: out <= 12'h000;
      20'h00ac3: out <= 12'h000;
      20'h00ac4: out <= 12'h000;
      20'h00ac5: out <= 12'h000;
      20'h00ac6: out <= 12'h000;
      20'h00ac7: out <= 12'h000;
      20'h00ac8: out <= 12'h000;
      20'h00ac9: out <= 12'h000;
      20'h00aca: out <= 12'h000;
      20'h00acb: out <= 12'h000;
      20'h00acc: out <= 12'h000;
      20'h00acd: out <= 12'h000;
      20'h00ace: out <= 12'h000;
      20'h00acf: out <= 12'h000;
      20'h00ad0: out <= 12'h000;
      20'h00ad1: out <= 12'h000;
      20'h00ad2: out <= 12'h000;
      20'h00ad3: out <= 12'h000;
      20'h00ad4: out <= 12'h000;
      20'h00ad5: out <= 12'h000;
      20'h00ad6: out <= 12'h000;
      20'h00ad7: out <= 12'h000;
      20'h00ad8: out <= 12'h000;
      20'h00ad9: out <= 12'h000;
      20'h00ada: out <= 12'h000;
      20'h00adb: out <= 12'h000;
      20'h00adc: out <= 12'h000;
      20'h00add: out <= 12'h000;
      20'h00ade: out <= 12'h000;
      20'h00adf: out <= 12'h000;
      20'h00ae0: out <= 12'h000;
      20'h00ae1: out <= 12'h000;
      20'h00ae2: out <= 12'h000;
      20'h00ae3: out <= 12'h000;
      20'h00ae4: out <= 12'h000;
      20'h00ae5: out <= 12'h000;
      20'h00ae6: out <= 12'h000;
      20'h00ae7: out <= 12'h000;
      20'h00ae8: out <= 12'h000;
      20'h00ae9: out <= 12'h000;
      20'h00aea: out <= 12'h000;
      20'h00aeb: out <= 12'h000;
      20'h00aec: out <= 12'h000;
      20'h00aed: out <= 12'h000;
      20'h00aee: out <= 12'h000;
      20'h00aef: out <= 12'h000;
      20'h00af0: out <= 12'h222;
      20'h00af1: out <= 12'h222;
      20'h00af2: out <= 12'h16d;
      20'h00af3: out <= 12'hfff;
      20'h00af4: out <= 12'h6af;
      20'h00af5: out <= 12'h6af;
      20'h00af6: out <= 12'h16d;
      20'h00af7: out <= 12'h16d;
      20'h00af8: out <= 12'h16d;
      20'h00af9: out <= 12'h6af;
      20'h00afa: out <= 12'hfff;
      20'h00afb: out <= 12'h16d;
      20'h00afc: out <= 12'h222;
      20'h00afd: out <= 12'h222;
      20'h00afe: out <= 12'h222;
      20'h00aff: out <= 12'h222;
      20'h00b00: out <= 12'h000;
      20'h00b01: out <= 12'h000;
      20'h00b02: out <= 12'h16d;
      20'h00b03: out <= 12'hfff;
      20'h00b04: out <= 12'h6af;
      20'h00b05: out <= 12'h6af;
      20'h00b06: out <= 12'h16d;
      20'h00b07: out <= 12'h16d;
      20'h00b08: out <= 12'h16d;
      20'h00b09: out <= 12'h6af;
      20'h00b0a: out <= 12'hfff;
      20'h00b0b: out <= 12'h16d;
      20'h00b0c: out <= 12'h000;
      20'h00b0d: out <= 12'h000;
      20'h00b0e: out <= 12'h000;
      20'h00b0f: out <= 12'h000;
      20'h00b10: out <= 12'h222;
      20'h00b11: out <= 12'h6af;
      20'h00b12: out <= 12'hfff;
      20'h00b13: out <= 12'h16d;
      20'h00b14: out <= 12'h6af;
      20'h00b15: out <= 12'h6af;
      20'h00b16: out <= 12'h16d;
      20'h00b17: out <= 12'h16d;
      20'h00b18: out <= 12'h6af;
      20'h00b19: out <= 12'h16d;
      20'h00b1a: out <= 12'h16d;
      20'h00b1b: out <= 12'h6af;
      20'h00b1c: out <= 12'h6af;
      20'h00b1d: out <= 12'h16d;
      20'h00b1e: out <= 12'hfff;
      20'h00b1f: out <= 12'h6af;
      20'h00b20: out <= 12'h000;
      20'h00b21: out <= 12'h6af;
      20'h00b22: out <= 12'h16d;
      20'h00b23: out <= 12'h16d;
      20'h00b24: out <= 12'h6af;
      20'h00b25: out <= 12'h6af;
      20'h00b26: out <= 12'h16d;
      20'h00b27: out <= 12'h16d;
      20'h00b28: out <= 12'h6af;
      20'h00b29: out <= 12'h16d;
      20'h00b2a: out <= 12'h16d;
      20'h00b2b: out <= 12'h6af;
      20'h00b2c: out <= 12'h6af;
      20'h00b2d: out <= 12'h16d;
      20'h00b2e: out <= 12'h16d;
      20'h00b2f: out <= 12'h6af;
      20'h00b30: out <= 12'h222;
      20'h00b31: out <= 12'h222;
      20'h00b32: out <= 12'h222;
      20'h00b33: out <= 12'h222;
      20'h00b34: out <= 12'h16d;
      20'h00b35: out <= 12'hfff;
      20'h00b36: out <= 12'h6af;
      20'h00b37: out <= 12'h16d;
      20'h00b38: out <= 12'h16d;
      20'h00b39: out <= 12'h16d;
      20'h00b3a: out <= 12'h6af;
      20'h00b3b: out <= 12'h6af;
      20'h00b3c: out <= 12'hfff;
      20'h00b3d: out <= 12'h16d;
      20'h00b3e: out <= 12'h222;
      20'h00b3f: out <= 12'h222;
      20'h00b40: out <= 12'h000;
      20'h00b41: out <= 12'h000;
      20'h00b42: out <= 12'h000;
      20'h00b43: out <= 12'h000;
      20'h00b44: out <= 12'h16d;
      20'h00b45: out <= 12'hfff;
      20'h00b46: out <= 12'h6af;
      20'h00b47: out <= 12'h16d;
      20'h00b48: out <= 12'h16d;
      20'h00b49: out <= 12'h16d;
      20'h00b4a: out <= 12'h6af;
      20'h00b4b: out <= 12'h6af;
      20'h00b4c: out <= 12'hfff;
      20'h00b4d: out <= 12'h16d;
      20'h00b4e: out <= 12'h000;
      20'h00b4f: out <= 12'h000;
      20'h00b50: out <= 12'h222;
      20'h00b51: out <= 12'h6af;
      20'h00b52: out <= 12'h16d;
      20'h00b53: out <= 12'h16d;
      20'h00b54: out <= 12'h16d;
      20'h00b55: out <= 12'hfff;
      20'h00b56: out <= 12'h6af;
      20'h00b57: out <= 12'h16d;
      20'h00b58: out <= 12'h16d;
      20'h00b59: out <= 12'h16d;
      20'h00b5a: out <= 12'h6af;
      20'h00b5b: out <= 12'hfff;
      20'h00b5c: out <= 12'h16d;
      20'h00b5d: out <= 12'h16d;
      20'h00b5e: out <= 12'h16d;
      20'h00b5f: out <= 12'h6af;
      20'h00b60: out <= 12'h000;
      20'h00b61: out <= 12'h6af;
      20'h00b62: out <= 12'hfff;
      20'h00b63: out <= 12'h16d;
      20'h00b64: out <= 12'h16d;
      20'h00b65: out <= 12'hfff;
      20'h00b66: out <= 12'h6af;
      20'h00b67: out <= 12'h16d;
      20'h00b68: out <= 12'h16d;
      20'h00b69: out <= 12'h16d;
      20'h00b6a: out <= 12'h6af;
      20'h00b6b: out <= 12'hfff;
      20'h00b6c: out <= 12'h16d;
      20'h00b6d: out <= 12'h16d;
      20'h00b6e: out <= 12'hfff;
      20'h00b6f: out <= 12'h6af;
      20'h00b70: out <= 12'h603;
      20'h00b71: out <= 12'h603;
      20'h00b72: out <= 12'h603;
      20'h00b73: out <= 12'h603;
      20'h00b74: out <= 12'hf87;
      20'h00b75: out <= 12'hf87;
      20'h00b76: out <= 12'hf87;
      20'h00b77: out <= 12'hee9;
      20'h00b78: out <= 12'hb27;
      20'h00b79: out <= 12'hf87;
      20'h00b7a: out <= 12'hf87;
      20'h00b7b: out <= 12'hf87;
      20'h00b7c: out <= 12'hf87;
      20'h00b7d: out <= 12'hf87;
      20'h00b7e: out <= 12'hf87;
      20'h00b7f: out <= 12'hee9;
      20'h00b80: out <= 12'hb27;
      20'h00b81: out <= 12'hf87;
      20'h00b82: out <= 12'hf87;
      20'h00b83: out <= 12'hf87;
      20'h00b84: out <= 12'h000;
      20'h00b85: out <= 12'h000;
      20'h00b86: out <= 12'h000;
      20'h00b87: out <= 12'h000;
      20'h00b88: out <= 12'h000;
      20'h00b89: out <= 12'h000;
      20'h00b8a: out <= 12'h000;
      20'h00b8b: out <= 12'h000;
      20'h00b8c: out <= 12'hf87;
      20'h00b8d: out <= 12'hf87;
      20'h00b8e: out <= 12'hf87;
      20'h00b8f: out <= 12'hee9;
      20'h00b90: out <= 12'hb27;
      20'h00b91: out <= 12'hf87;
      20'h00b92: out <= 12'hf87;
      20'h00b93: out <= 12'hf87;
      20'h00b94: out <= 12'hf87;
      20'h00b95: out <= 12'hf87;
      20'h00b96: out <= 12'hf87;
      20'h00b97: out <= 12'hee9;
      20'h00b98: out <= 12'hb27;
      20'h00b99: out <= 12'hf87;
      20'h00b9a: out <= 12'hf87;
      20'h00b9b: out <= 12'hf87;
      20'h00b9c: out <= 12'hf87;
      20'h00b9d: out <= 12'hf87;
      20'h00b9e: out <= 12'hf87;
      20'h00b9f: out <= 12'hee9;
      20'h00ba0: out <= 12'hb27;
      20'h00ba1: out <= 12'hf87;
      20'h00ba2: out <= 12'hf87;
      20'h00ba3: out <= 12'hf87;
      20'h00ba4: out <= 12'hf87;
      20'h00ba5: out <= 12'hf87;
      20'h00ba6: out <= 12'hf87;
      20'h00ba7: out <= 12'hee9;
      20'h00ba8: out <= 12'hb27;
      20'h00ba9: out <= 12'hf87;
      20'h00baa: out <= 12'hf87;
      20'h00bab: out <= 12'hf87;
      20'h00bac: out <= 12'h000;
      20'h00bad: out <= 12'h000;
      20'h00bae: out <= 12'h000;
      20'h00baf: out <= 12'h000;
      20'h00bb0: out <= 12'h000;
      20'h00bb1: out <= 12'h000;
      20'h00bb2: out <= 12'h000;
      20'h00bb3: out <= 12'h000;
      20'h00bb4: out <= 12'h000;
      20'h00bb5: out <= 12'h000;
      20'h00bb6: out <= 12'h000;
      20'h00bb7: out <= 12'h000;
      20'h00bb8: out <= 12'h000;
      20'h00bb9: out <= 12'h000;
      20'h00bba: out <= 12'h000;
      20'h00bbb: out <= 12'h000;
      20'h00bbc: out <= 12'h000;
      20'h00bbd: out <= 12'h000;
      20'h00bbe: out <= 12'h000;
      20'h00bbf: out <= 12'h000;
      20'h00bc0: out <= 12'h000;
      20'h00bc1: out <= 12'h000;
      20'h00bc2: out <= 12'h000;
      20'h00bc3: out <= 12'h000;
      20'h00bc4: out <= 12'h603;
      20'h00bc5: out <= 12'h603;
      20'h00bc6: out <= 12'h603;
      20'h00bc7: out <= 12'h603;
      20'h00bc8: out <= 12'hee9;
      20'h00bc9: out <= 12'hf87;
      20'h00bca: out <= 12'hee9;
      20'h00bcb: out <= 12'hee9;
      20'h00bcc: out <= 12'hee9;
      20'h00bcd: out <= 12'hb27;
      20'h00bce: out <= 12'hf87;
      20'h00bcf: out <= 12'hb27;
      20'h00bd0: out <= 12'h000;
      20'h00bd1: out <= 12'h000;
      20'h00bd2: out <= 12'h000;
      20'h00bd3: out <= 12'h000;
      20'h00bd4: out <= 12'h000;
      20'h00bd5: out <= 12'h000;
      20'h00bd6: out <= 12'h000;
      20'h00bd7: out <= 12'h000;
      20'h00bd8: out <= 12'h000;
      20'h00bd9: out <= 12'h000;
      20'h00bda: out <= 12'h000;
      20'h00bdb: out <= 12'h000;
      20'h00bdc: out <= 12'h000;
      20'h00bdd: out <= 12'h000;
      20'h00bde: out <= 12'h000;
      20'h00bdf: out <= 12'h000;
      20'h00be0: out <= 12'h000;
      20'h00be1: out <= 12'h000;
      20'h00be2: out <= 12'h000;
      20'h00be3: out <= 12'h000;
      20'h00be4: out <= 12'h000;
      20'h00be5: out <= 12'h000;
      20'h00be6: out <= 12'h000;
      20'h00be7: out <= 12'h000;
      20'h00be8: out <= 12'h000;
      20'h00be9: out <= 12'h000;
      20'h00bea: out <= 12'h000;
      20'h00beb: out <= 12'h000;
      20'h00bec: out <= 12'h000;
      20'h00bed: out <= 12'h000;
      20'h00bee: out <= 12'h000;
      20'h00bef: out <= 12'h000;
      20'h00bf0: out <= 12'h000;
      20'h00bf1: out <= 12'h000;
      20'h00bf2: out <= 12'h000;
      20'h00bf3: out <= 12'h000;
      20'h00bf4: out <= 12'h000;
      20'h00bf5: out <= 12'h000;
      20'h00bf6: out <= 12'h000;
      20'h00bf7: out <= 12'h000;
      20'h00bf8: out <= 12'h000;
      20'h00bf9: out <= 12'h000;
      20'h00bfa: out <= 12'h000;
      20'h00bfb: out <= 12'h000;
      20'h00bfc: out <= 12'h000;
      20'h00bfd: out <= 12'h000;
      20'h00bfe: out <= 12'h000;
      20'h00bff: out <= 12'h000;
      20'h00c00: out <= 12'h000;
      20'h00c01: out <= 12'h000;
      20'h00c02: out <= 12'h000;
      20'h00c03: out <= 12'h000;
      20'h00c04: out <= 12'h000;
      20'h00c05: out <= 12'h000;
      20'h00c06: out <= 12'h000;
      20'h00c07: out <= 12'h000;
      20'h00c08: out <= 12'h222;
      20'h00c09: out <= 12'h222;
      20'h00c0a: out <= 12'h222;
      20'h00c0b: out <= 12'h16d;
      20'h00c0c: out <= 12'hfff;
      20'h00c0d: out <= 12'h6af;
      20'h00c0e: out <= 12'h6af;
      20'h00c0f: out <= 12'h6af;
      20'h00c10: out <= 12'h6af;
      20'h00c11: out <= 12'hfff;
      20'h00c12: out <= 12'h16d;
      20'h00c13: out <= 12'h222;
      20'h00c14: out <= 12'h222;
      20'h00c15: out <= 12'h222;
      20'h00c16: out <= 12'h222;
      20'h00c17: out <= 12'h222;
      20'h00c18: out <= 12'h000;
      20'h00c19: out <= 12'h000;
      20'h00c1a: out <= 12'h000;
      20'h00c1b: out <= 12'h16d;
      20'h00c1c: out <= 12'hfff;
      20'h00c1d: out <= 12'h6af;
      20'h00c1e: out <= 12'h6af;
      20'h00c1f: out <= 12'h6af;
      20'h00c20: out <= 12'h6af;
      20'h00c21: out <= 12'hfff;
      20'h00c22: out <= 12'h16d;
      20'h00c23: out <= 12'h000;
      20'h00c24: out <= 12'h000;
      20'h00c25: out <= 12'h000;
      20'h00c26: out <= 12'h000;
      20'h00c27: out <= 12'h000;
      20'h00c28: out <= 12'h222;
      20'h00c29: out <= 12'h6af;
      20'h00c2a: out <= 12'h16d;
      20'h00c2b: out <= 12'h16d;
      20'h00c2c: out <= 12'hfff;
      20'h00c2d: out <= 12'h6af;
      20'h00c2e: out <= 12'h6af;
      20'h00c2f: out <= 12'h16d;
      20'h00c30: out <= 12'h16d;
      20'h00c31: out <= 12'h16d;
      20'h00c32: out <= 12'h6af;
      20'h00c33: out <= 12'h6af;
      20'h00c34: out <= 12'hfff;
      20'h00c35: out <= 12'h16d;
      20'h00c36: out <= 12'h16d;
      20'h00c37: out <= 12'h6af;
      20'h00c38: out <= 12'h000;
      20'h00c39: out <= 12'h6af;
      20'h00c3a: out <= 12'hfff;
      20'h00c3b: out <= 12'h16d;
      20'h00c3c: out <= 12'hfff;
      20'h00c3d: out <= 12'h6af;
      20'h00c3e: out <= 12'h6af;
      20'h00c3f: out <= 12'h16d;
      20'h00c40: out <= 12'h16d;
      20'h00c41: out <= 12'h16d;
      20'h00c42: out <= 12'h6af;
      20'h00c43: out <= 12'h6af;
      20'h00c44: out <= 12'hfff;
      20'h00c45: out <= 12'h16d;
      20'h00c46: out <= 12'hfff;
      20'h00c47: out <= 12'h6af;
      20'h00c48: out <= 12'h222;
      20'h00c49: out <= 12'h222;
      20'h00c4a: out <= 12'h222;
      20'h00c4b: out <= 12'h222;
      20'h00c4c: out <= 12'h222;
      20'h00c4d: out <= 12'h16d;
      20'h00c4e: out <= 12'hfff;
      20'h00c4f: out <= 12'h6af;
      20'h00c50: out <= 12'h6af;
      20'h00c51: out <= 12'h6af;
      20'h00c52: out <= 12'h6af;
      20'h00c53: out <= 12'hfff;
      20'h00c54: out <= 12'h16d;
      20'h00c55: out <= 12'h222;
      20'h00c56: out <= 12'h222;
      20'h00c57: out <= 12'h222;
      20'h00c58: out <= 12'h000;
      20'h00c59: out <= 12'h000;
      20'h00c5a: out <= 12'h000;
      20'h00c5b: out <= 12'h000;
      20'h00c5c: out <= 12'h000;
      20'h00c5d: out <= 12'h16d;
      20'h00c5e: out <= 12'hfff;
      20'h00c5f: out <= 12'h6af;
      20'h00c60: out <= 12'h6af;
      20'h00c61: out <= 12'h6af;
      20'h00c62: out <= 12'h6af;
      20'h00c63: out <= 12'hfff;
      20'h00c64: out <= 12'h16d;
      20'h00c65: out <= 12'h000;
      20'h00c66: out <= 12'h000;
      20'h00c67: out <= 12'h000;
      20'h00c68: out <= 12'h222;
      20'h00c69: out <= 12'h6af;
      20'h00c6a: out <= 12'hfff;
      20'h00c6b: out <= 12'h6af;
      20'h00c6c: out <= 12'h222;
      20'h00c6d: out <= 12'h16d;
      20'h00c6e: out <= 12'h16d;
      20'h00c6f: out <= 12'h16d;
      20'h00c70: out <= 12'hfff;
      20'h00c71: out <= 12'h16d;
      20'h00c72: out <= 12'h16d;
      20'h00c73: out <= 12'h16d;
      20'h00c74: out <= 12'h222;
      20'h00c75: out <= 12'h6af;
      20'h00c76: out <= 12'hfff;
      20'h00c77: out <= 12'h6af;
      20'h00c78: out <= 12'h000;
      20'h00c79: out <= 12'h6af;
      20'h00c7a: out <= 12'h16d;
      20'h00c7b: out <= 12'h6af;
      20'h00c7c: out <= 12'h000;
      20'h00c7d: out <= 12'h16d;
      20'h00c7e: out <= 12'h16d;
      20'h00c7f: out <= 12'h16d;
      20'h00c80: out <= 12'hfff;
      20'h00c81: out <= 12'h16d;
      20'h00c82: out <= 12'h16d;
      20'h00c83: out <= 12'h16d;
      20'h00c84: out <= 12'h000;
      20'h00c85: out <= 12'h6af;
      20'h00c86: out <= 12'h16d;
      20'h00c87: out <= 12'h6af;
      20'h00c88: out <= 12'h603;
      20'h00c89: out <= 12'h603;
      20'h00c8a: out <= 12'h603;
      20'h00c8b: out <= 12'h603;
      20'h00c8c: out <= 12'hb27;
      20'h00c8d: out <= 12'hb27;
      20'h00c8e: out <= 12'hb27;
      20'h00c8f: out <= 12'hb27;
      20'h00c90: out <= 12'hb27;
      20'h00c91: out <= 12'hb27;
      20'h00c92: out <= 12'hb27;
      20'h00c93: out <= 12'hb27;
      20'h00c94: out <= 12'hb27;
      20'h00c95: out <= 12'hb27;
      20'h00c96: out <= 12'hb27;
      20'h00c97: out <= 12'hb27;
      20'h00c98: out <= 12'hb27;
      20'h00c99: out <= 12'hb27;
      20'h00c9a: out <= 12'hb27;
      20'h00c9b: out <= 12'hb27;
      20'h00c9c: out <= 12'h000;
      20'h00c9d: out <= 12'h000;
      20'h00c9e: out <= 12'h000;
      20'h00c9f: out <= 12'h000;
      20'h00ca0: out <= 12'h000;
      20'h00ca1: out <= 12'h000;
      20'h00ca2: out <= 12'h000;
      20'h00ca3: out <= 12'h000;
      20'h00ca4: out <= 12'hb27;
      20'h00ca5: out <= 12'hb27;
      20'h00ca6: out <= 12'hb27;
      20'h00ca7: out <= 12'hb27;
      20'h00ca8: out <= 12'hb27;
      20'h00ca9: out <= 12'hb27;
      20'h00caa: out <= 12'hb27;
      20'h00cab: out <= 12'hb27;
      20'h00cac: out <= 12'hb27;
      20'h00cad: out <= 12'hb27;
      20'h00cae: out <= 12'hb27;
      20'h00caf: out <= 12'hb27;
      20'h00cb0: out <= 12'hb27;
      20'h00cb1: out <= 12'hb27;
      20'h00cb2: out <= 12'hb27;
      20'h00cb3: out <= 12'hb27;
      20'h00cb4: out <= 12'hb27;
      20'h00cb5: out <= 12'hb27;
      20'h00cb6: out <= 12'hb27;
      20'h00cb7: out <= 12'hb27;
      20'h00cb8: out <= 12'hb27;
      20'h00cb9: out <= 12'hb27;
      20'h00cba: out <= 12'hb27;
      20'h00cbb: out <= 12'hb27;
      20'h00cbc: out <= 12'hb27;
      20'h00cbd: out <= 12'hb27;
      20'h00cbe: out <= 12'hb27;
      20'h00cbf: out <= 12'hb27;
      20'h00cc0: out <= 12'hb27;
      20'h00cc1: out <= 12'hb27;
      20'h00cc2: out <= 12'hb27;
      20'h00cc3: out <= 12'hb27;
      20'h00cc4: out <= 12'h000;
      20'h00cc5: out <= 12'h000;
      20'h00cc6: out <= 12'h000;
      20'h00cc7: out <= 12'h000;
      20'h00cc8: out <= 12'h000;
      20'h00cc9: out <= 12'h000;
      20'h00cca: out <= 12'h000;
      20'h00ccb: out <= 12'h000;
      20'h00ccc: out <= 12'h000;
      20'h00ccd: out <= 12'h000;
      20'h00cce: out <= 12'h000;
      20'h00ccf: out <= 12'h000;
      20'h00cd0: out <= 12'h000;
      20'h00cd1: out <= 12'h000;
      20'h00cd2: out <= 12'h000;
      20'h00cd3: out <= 12'h000;
      20'h00cd4: out <= 12'h000;
      20'h00cd5: out <= 12'h000;
      20'h00cd6: out <= 12'h000;
      20'h00cd7: out <= 12'h000;
      20'h00cd8: out <= 12'h000;
      20'h00cd9: out <= 12'h000;
      20'h00cda: out <= 12'h000;
      20'h00cdb: out <= 12'h000;
      20'h00cdc: out <= 12'h603;
      20'h00cdd: out <= 12'h603;
      20'h00cde: out <= 12'h603;
      20'h00cdf: out <= 12'h603;
      20'h00ce0: out <= 12'hee9;
      20'h00ce1: out <= 12'hf87;
      20'h00ce2: out <= 12'hee9;
      20'h00ce3: out <= 12'hf87;
      20'h00ce4: out <= 12'hf87;
      20'h00ce5: out <= 12'hb27;
      20'h00ce6: out <= 12'hf87;
      20'h00ce7: out <= 12'hb27;
      20'h00ce8: out <= 12'h000;
      20'h00ce9: out <= 12'h000;
      20'h00cea: out <= 12'h000;
      20'h00ceb: out <= 12'h000;
      20'h00cec: out <= 12'h000;
      20'h00ced: out <= 12'h000;
      20'h00cee: out <= 12'h000;
      20'h00cef: out <= 12'h000;
      20'h00cf0: out <= 12'h000;
      20'h00cf1: out <= 12'h000;
      20'h00cf2: out <= 12'h000;
      20'h00cf3: out <= 12'h000;
      20'h00cf4: out <= 12'h000;
      20'h00cf5: out <= 12'h000;
      20'h00cf6: out <= 12'h000;
      20'h00cf7: out <= 12'h000;
      20'h00cf8: out <= 12'h000;
      20'h00cf9: out <= 12'h000;
      20'h00cfa: out <= 12'h000;
      20'h00cfb: out <= 12'h000;
      20'h00cfc: out <= 12'h000;
      20'h00cfd: out <= 12'h000;
      20'h00cfe: out <= 12'h000;
      20'h00cff: out <= 12'h000;
      20'h00d00: out <= 12'h000;
      20'h00d01: out <= 12'h000;
      20'h00d02: out <= 12'h000;
      20'h00d03: out <= 12'h000;
      20'h00d04: out <= 12'h000;
      20'h00d05: out <= 12'h000;
      20'h00d06: out <= 12'h000;
      20'h00d07: out <= 12'h000;
      20'h00d08: out <= 12'h000;
      20'h00d09: out <= 12'h000;
      20'h00d0a: out <= 12'h000;
      20'h00d0b: out <= 12'h000;
      20'h00d0c: out <= 12'h000;
      20'h00d0d: out <= 12'h000;
      20'h00d0e: out <= 12'h000;
      20'h00d0f: out <= 12'h000;
      20'h00d10: out <= 12'h000;
      20'h00d11: out <= 12'h000;
      20'h00d12: out <= 12'h000;
      20'h00d13: out <= 12'h000;
      20'h00d14: out <= 12'h000;
      20'h00d15: out <= 12'h000;
      20'h00d16: out <= 12'h000;
      20'h00d17: out <= 12'h000;
      20'h00d18: out <= 12'h000;
      20'h00d19: out <= 12'h000;
      20'h00d1a: out <= 12'h000;
      20'h00d1b: out <= 12'h000;
      20'h00d1c: out <= 12'h000;
      20'h00d1d: out <= 12'h000;
      20'h00d1e: out <= 12'h000;
      20'h00d1f: out <= 12'h000;
      20'h00d20: out <= 12'h222;
      20'h00d21: out <= 12'h6af;
      20'h00d22: out <= 12'h6af;
      20'h00d23: out <= 12'h6af;
      20'h00d24: out <= 12'h16d;
      20'h00d25: out <= 12'h16d;
      20'h00d26: out <= 12'h16d;
      20'h00d27: out <= 12'h16d;
      20'h00d28: out <= 12'h16d;
      20'h00d29: out <= 12'h16d;
      20'h00d2a: out <= 12'h16d;
      20'h00d2b: out <= 12'h6af;
      20'h00d2c: out <= 12'h6af;
      20'h00d2d: out <= 12'h222;
      20'h00d2e: out <= 12'h222;
      20'h00d2f: out <= 12'h222;
      20'h00d30: out <= 12'h000;
      20'h00d31: out <= 12'h6af;
      20'h00d32: out <= 12'h6af;
      20'h00d33: out <= 12'h6af;
      20'h00d34: out <= 12'h16d;
      20'h00d35: out <= 12'h16d;
      20'h00d36: out <= 12'h16d;
      20'h00d37: out <= 12'h16d;
      20'h00d38: out <= 12'h16d;
      20'h00d39: out <= 12'h16d;
      20'h00d3a: out <= 12'h16d;
      20'h00d3b: out <= 12'h6af;
      20'h00d3c: out <= 12'h6af;
      20'h00d3d: out <= 12'h000;
      20'h00d3e: out <= 12'h000;
      20'h00d3f: out <= 12'h000;
      20'h00d40: out <= 12'h222;
      20'h00d41: out <= 12'h6af;
      20'h00d42: out <= 12'hfff;
      20'h00d43: out <= 12'h6af;
      20'h00d44: out <= 12'h16d;
      20'h00d45: out <= 12'hfff;
      20'h00d46: out <= 12'h6af;
      20'h00d47: out <= 12'h6af;
      20'h00d48: out <= 12'h6af;
      20'h00d49: out <= 12'h6af;
      20'h00d4a: out <= 12'h6af;
      20'h00d4b: out <= 12'hfff;
      20'h00d4c: out <= 12'h16d;
      20'h00d4d: out <= 12'h6af;
      20'h00d4e: out <= 12'hfff;
      20'h00d4f: out <= 12'h6af;
      20'h00d50: out <= 12'h000;
      20'h00d51: out <= 12'h6af;
      20'h00d52: out <= 12'h16d;
      20'h00d53: out <= 12'h6af;
      20'h00d54: out <= 12'h16d;
      20'h00d55: out <= 12'hfff;
      20'h00d56: out <= 12'h6af;
      20'h00d57: out <= 12'h6af;
      20'h00d58: out <= 12'h6af;
      20'h00d59: out <= 12'h6af;
      20'h00d5a: out <= 12'h6af;
      20'h00d5b: out <= 12'hfff;
      20'h00d5c: out <= 12'h16d;
      20'h00d5d: out <= 12'h6af;
      20'h00d5e: out <= 12'h16d;
      20'h00d5f: out <= 12'h6af;
      20'h00d60: out <= 12'h222;
      20'h00d61: out <= 12'h222;
      20'h00d62: out <= 12'h222;
      20'h00d63: out <= 12'h6af;
      20'h00d64: out <= 12'h6af;
      20'h00d65: out <= 12'h16d;
      20'h00d66: out <= 12'h16d;
      20'h00d67: out <= 12'h16d;
      20'h00d68: out <= 12'h16d;
      20'h00d69: out <= 12'h16d;
      20'h00d6a: out <= 12'h16d;
      20'h00d6b: out <= 12'h16d;
      20'h00d6c: out <= 12'h6af;
      20'h00d6d: out <= 12'h6af;
      20'h00d6e: out <= 12'h6af;
      20'h00d6f: out <= 12'h222;
      20'h00d70: out <= 12'h000;
      20'h00d71: out <= 12'h000;
      20'h00d72: out <= 12'h000;
      20'h00d73: out <= 12'h6af;
      20'h00d74: out <= 12'h6af;
      20'h00d75: out <= 12'h16d;
      20'h00d76: out <= 12'h16d;
      20'h00d77: out <= 12'h16d;
      20'h00d78: out <= 12'h16d;
      20'h00d79: out <= 12'h16d;
      20'h00d7a: out <= 12'h16d;
      20'h00d7b: out <= 12'h16d;
      20'h00d7c: out <= 12'h6af;
      20'h00d7d: out <= 12'h6af;
      20'h00d7e: out <= 12'h6af;
      20'h00d7f: out <= 12'h000;
      20'h00d80: out <= 12'h222;
      20'h00d81: out <= 12'h6af;
      20'h00d82: out <= 12'h16d;
      20'h00d83: out <= 12'h6af;
      20'h00d84: out <= 12'h222;
      20'h00d85: out <= 12'h222;
      20'h00d86: out <= 12'h222;
      20'h00d87: out <= 12'h16d;
      20'h00d88: out <= 12'hfff;
      20'h00d89: out <= 12'h16d;
      20'h00d8a: out <= 12'h222;
      20'h00d8b: out <= 12'h222;
      20'h00d8c: out <= 12'h222;
      20'h00d8d: out <= 12'h6af;
      20'h00d8e: out <= 12'h16d;
      20'h00d8f: out <= 12'h6af;
      20'h00d90: out <= 12'h000;
      20'h00d91: out <= 12'h6af;
      20'h00d92: out <= 12'hfff;
      20'h00d93: out <= 12'h6af;
      20'h00d94: out <= 12'h000;
      20'h00d95: out <= 12'h000;
      20'h00d96: out <= 12'h000;
      20'h00d97: out <= 12'h16d;
      20'h00d98: out <= 12'hfff;
      20'h00d99: out <= 12'h16d;
      20'h00d9a: out <= 12'h000;
      20'h00d9b: out <= 12'h000;
      20'h00d9c: out <= 12'h000;
      20'h00d9d: out <= 12'h6af;
      20'h00d9e: out <= 12'hfff;
      20'h00d9f: out <= 12'h6af;
      20'h00da0: out <= 12'h603;
      20'h00da1: out <= 12'h603;
      20'h00da2: out <= 12'h603;
      20'h00da3: out <= 12'h603;
      20'h00da4: out <= 12'hb27;
      20'h00da5: out <= 12'hee9;
      20'h00da6: out <= 12'hee9;
      20'h00da7: out <= 12'hee9;
      20'h00da8: out <= 12'hee9;
      20'h00da9: out <= 12'hee9;
      20'h00daa: out <= 12'hee9;
      20'h00dab: out <= 12'hee9;
      20'h00dac: out <= 12'hb27;
      20'h00dad: out <= 12'hee9;
      20'h00dae: out <= 12'hee9;
      20'h00daf: out <= 12'hee9;
      20'h00db0: out <= 12'hee9;
      20'h00db1: out <= 12'hee9;
      20'h00db2: out <= 12'hee9;
      20'h00db3: out <= 12'hee9;
      20'h00db4: out <= 12'h000;
      20'h00db5: out <= 12'h000;
      20'h00db6: out <= 12'h000;
      20'h00db7: out <= 12'h000;
      20'h00db8: out <= 12'h000;
      20'h00db9: out <= 12'h000;
      20'h00dba: out <= 12'h000;
      20'h00dbb: out <= 12'h000;
      20'h00dbc: out <= 12'hb27;
      20'h00dbd: out <= 12'hee9;
      20'h00dbe: out <= 12'hee9;
      20'h00dbf: out <= 12'hee9;
      20'h00dc0: out <= 12'hee9;
      20'h00dc1: out <= 12'hee9;
      20'h00dc2: out <= 12'hee9;
      20'h00dc3: out <= 12'hee9;
      20'h00dc4: out <= 12'hb27;
      20'h00dc5: out <= 12'hee9;
      20'h00dc6: out <= 12'hee9;
      20'h00dc7: out <= 12'hee9;
      20'h00dc8: out <= 12'hee9;
      20'h00dc9: out <= 12'hee9;
      20'h00dca: out <= 12'hee9;
      20'h00dcb: out <= 12'hee9;
      20'h00dcc: out <= 12'hb27;
      20'h00dcd: out <= 12'hee9;
      20'h00dce: out <= 12'hee9;
      20'h00dcf: out <= 12'hee9;
      20'h00dd0: out <= 12'hee9;
      20'h00dd1: out <= 12'hee9;
      20'h00dd2: out <= 12'hee9;
      20'h00dd3: out <= 12'hee9;
      20'h00dd4: out <= 12'hb27;
      20'h00dd5: out <= 12'hee9;
      20'h00dd6: out <= 12'hee9;
      20'h00dd7: out <= 12'hee9;
      20'h00dd8: out <= 12'hee9;
      20'h00dd9: out <= 12'hee9;
      20'h00dda: out <= 12'hee9;
      20'h00ddb: out <= 12'hee9;
      20'h00ddc: out <= 12'h000;
      20'h00ddd: out <= 12'h000;
      20'h00dde: out <= 12'h000;
      20'h00ddf: out <= 12'h000;
      20'h00de0: out <= 12'h000;
      20'h00de1: out <= 12'h000;
      20'h00de2: out <= 12'h000;
      20'h00de3: out <= 12'h000;
      20'h00de4: out <= 12'h000;
      20'h00de5: out <= 12'h000;
      20'h00de6: out <= 12'h000;
      20'h00de7: out <= 12'h000;
      20'h00de8: out <= 12'h000;
      20'h00de9: out <= 12'h000;
      20'h00dea: out <= 12'h000;
      20'h00deb: out <= 12'h000;
      20'h00dec: out <= 12'h000;
      20'h00ded: out <= 12'h000;
      20'h00dee: out <= 12'h000;
      20'h00def: out <= 12'h000;
      20'h00df0: out <= 12'h000;
      20'h00df1: out <= 12'h000;
      20'h00df2: out <= 12'h000;
      20'h00df3: out <= 12'h000;
      20'h00df4: out <= 12'h603;
      20'h00df5: out <= 12'h603;
      20'h00df6: out <= 12'h603;
      20'h00df7: out <= 12'h603;
      20'h00df8: out <= 12'hee9;
      20'h00df9: out <= 12'hf87;
      20'h00dfa: out <= 12'hee9;
      20'h00dfb: out <= 12'hf87;
      20'h00dfc: out <= 12'hf87;
      20'h00dfd: out <= 12'hb27;
      20'h00dfe: out <= 12'hf87;
      20'h00dff: out <= 12'hb27;
      20'h00e00: out <= 12'h000;
      20'h00e01: out <= 12'h000;
      20'h00e02: out <= 12'h000;
      20'h00e03: out <= 12'h000;
      20'h00e04: out <= 12'h000;
      20'h00e05: out <= 12'h000;
      20'h00e06: out <= 12'h000;
      20'h00e07: out <= 12'h000;
      20'h00e08: out <= 12'h000;
      20'h00e09: out <= 12'h000;
      20'h00e0a: out <= 12'h000;
      20'h00e0b: out <= 12'h000;
      20'h00e0c: out <= 12'h000;
      20'h00e0d: out <= 12'h000;
      20'h00e0e: out <= 12'h000;
      20'h00e0f: out <= 12'h000;
      20'h00e10: out <= 12'h000;
      20'h00e11: out <= 12'h000;
      20'h00e12: out <= 12'h000;
      20'h00e13: out <= 12'h000;
      20'h00e14: out <= 12'h000;
      20'h00e15: out <= 12'h000;
      20'h00e16: out <= 12'h000;
      20'h00e17: out <= 12'h000;
      20'h00e18: out <= 12'h000;
      20'h00e19: out <= 12'h000;
      20'h00e1a: out <= 12'h000;
      20'h00e1b: out <= 12'h000;
      20'h00e1c: out <= 12'h000;
      20'h00e1d: out <= 12'h000;
      20'h00e1e: out <= 12'h000;
      20'h00e1f: out <= 12'h000;
      20'h00e20: out <= 12'h000;
      20'h00e21: out <= 12'h000;
      20'h00e22: out <= 12'h000;
      20'h00e23: out <= 12'h000;
      20'h00e24: out <= 12'h000;
      20'h00e25: out <= 12'h000;
      20'h00e26: out <= 12'h000;
      20'h00e27: out <= 12'h000;
      20'h00e28: out <= 12'h000;
      20'h00e29: out <= 12'h000;
      20'h00e2a: out <= 12'h000;
      20'h00e2b: out <= 12'h000;
      20'h00e2c: out <= 12'h000;
      20'h00e2d: out <= 12'h000;
      20'h00e2e: out <= 12'h000;
      20'h00e2f: out <= 12'h000;
      20'h00e30: out <= 12'h000;
      20'h00e31: out <= 12'h000;
      20'h00e32: out <= 12'h000;
      20'h00e33: out <= 12'h000;
      20'h00e34: out <= 12'h000;
      20'h00e35: out <= 12'h000;
      20'h00e36: out <= 12'h000;
      20'h00e37: out <= 12'h000;
      20'h00e38: out <= 12'h222;
      20'h00e39: out <= 12'hfff;
      20'h00e3a: out <= 12'h16d;
      20'h00e3b: out <= 12'hfff;
      20'h00e3c: out <= 12'h16d;
      20'h00e3d: out <= 12'hfff;
      20'h00e3e: out <= 12'h16d;
      20'h00e3f: out <= 12'hfff;
      20'h00e40: out <= 12'h16d;
      20'h00e41: out <= 12'hfff;
      20'h00e42: out <= 12'h16d;
      20'h00e43: out <= 12'hfff;
      20'h00e44: out <= 12'h16d;
      20'h00e45: out <= 12'h222;
      20'h00e46: out <= 12'h222;
      20'h00e47: out <= 12'h222;
      20'h00e48: out <= 12'h000;
      20'h00e49: out <= 12'h6af;
      20'h00e4a: out <= 12'hfff;
      20'h00e4b: out <= 12'h16d;
      20'h00e4c: out <= 12'hfff;
      20'h00e4d: out <= 12'h16d;
      20'h00e4e: out <= 12'hfff;
      20'h00e4f: out <= 12'h16d;
      20'h00e50: out <= 12'hfff;
      20'h00e51: out <= 12'h16d;
      20'h00e52: out <= 12'hfff;
      20'h00e53: out <= 12'h16d;
      20'h00e54: out <= 12'hfff;
      20'h00e55: out <= 12'h000;
      20'h00e56: out <= 12'h000;
      20'h00e57: out <= 12'h000;
      20'h00e58: out <= 12'h222;
      20'h00e59: out <= 12'h6af;
      20'h00e5a: out <= 12'h16d;
      20'h00e5b: out <= 12'h6af;
      20'h00e5c: out <= 12'h222;
      20'h00e5d: out <= 12'h16d;
      20'h00e5e: out <= 12'h16d;
      20'h00e5f: out <= 12'h16d;
      20'h00e60: out <= 12'h16d;
      20'h00e61: out <= 12'h16d;
      20'h00e62: out <= 12'h16d;
      20'h00e63: out <= 12'h16d;
      20'h00e64: out <= 12'h222;
      20'h00e65: out <= 12'h6af;
      20'h00e66: out <= 12'h16d;
      20'h00e67: out <= 12'h6af;
      20'h00e68: out <= 12'h000;
      20'h00e69: out <= 12'h6af;
      20'h00e6a: out <= 12'hfff;
      20'h00e6b: out <= 12'h6af;
      20'h00e6c: out <= 12'h000;
      20'h00e6d: out <= 12'h16d;
      20'h00e6e: out <= 12'h16d;
      20'h00e6f: out <= 12'h16d;
      20'h00e70: out <= 12'h16d;
      20'h00e71: out <= 12'h16d;
      20'h00e72: out <= 12'h16d;
      20'h00e73: out <= 12'h16d;
      20'h00e74: out <= 12'h000;
      20'h00e75: out <= 12'h6af;
      20'h00e76: out <= 12'hfff;
      20'h00e77: out <= 12'h6af;
      20'h00e78: out <= 12'h222;
      20'h00e79: out <= 12'h222;
      20'h00e7a: out <= 12'h222;
      20'h00e7b: out <= 12'h16d;
      20'h00e7c: out <= 12'hfff;
      20'h00e7d: out <= 12'h16d;
      20'h00e7e: out <= 12'hfff;
      20'h00e7f: out <= 12'h16d;
      20'h00e80: out <= 12'hfff;
      20'h00e81: out <= 12'h16d;
      20'h00e82: out <= 12'hfff;
      20'h00e83: out <= 12'h16d;
      20'h00e84: out <= 12'hfff;
      20'h00e85: out <= 12'h16d;
      20'h00e86: out <= 12'hfff;
      20'h00e87: out <= 12'h222;
      20'h00e88: out <= 12'h000;
      20'h00e89: out <= 12'h000;
      20'h00e8a: out <= 12'h000;
      20'h00e8b: out <= 12'hfff;
      20'h00e8c: out <= 12'h16d;
      20'h00e8d: out <= 12'hfff;
      20'h00e8e: out <= 12'h16d;
      20'h00e8f: out <= 12'hfff;
      20'h00e90: out <= 12'h16d;
      20'h00e91: out <= 12'hfff;
      20'h00e92: out <= 12'h16d;
      20'h00e93: out <= 12'hfff;
      20'h00e94: out <= 12'h16d;
      20'h00e95: out <= 12'hfff;
      20'h00e96: out <= 12'h6af;
      20'h00e97: out <= 12'h000;
      20'h00e98: out <= 12'h222;
      20'h00e99: out <= 12'h222;
      20'h00e9a: out <= 12'h222;
      20'h00e9b: out <= 12'h222;
      20'h00e9c: out <= 12'h222;
      20'h00e9d: out <= 12'h222;
      20'h00e9e: out <= 12'h222;
      20'h00e9f: out <= 12'h16d;
      20'h00ea0: out <= 12'hfff;
      20'h00ea1: out <= 12'h16d;
      20'h00ea2: out <= 12'h222;
      20'h00ea3: out <= 12'h222;
      20'h00ea4: out <= 12'h222;
      20'h00ea5: out <= 12'h222;
      20'h00ea6: out <= 12'h222;
      20'h00ea7: out <= 12'h222;
      20'h00ea8: out <= 12'h000;
      20'h00ea9: out <= 12'h000;
      20'h00eaa: out <= 12'h000;
      20'h00eab: out <= 12'h000;
      20'h00eac: out <= 12'h000;
      20'h00ead: out <= 12'h000;
      20'h00eae: out <= 12'h000;
      20'h00eaf: out <= 12'h16d;
      20'h00eb0: out <= 12'hfff;
      20'h00eb1: out <= 12'h16d;
      20'h00eb2: out <= 12'h000;
      20'h00eb3: out <= 12'h000;
      20'h00eb4: out <= 12'h000;
      20'h00eb5: out <= 12'h000;
      20'h00eb6: out <= 12'h000;
      20'h00eb7: out <= 12'h000;
      20'h00eb8: out <= 12'h603;
      20'h00eb9: out <= 12'h603;
      20'h00eba: out <= 12'h603;
      20'h00ebb: out <= 12'h603;
      20'h00ebc: out <= 12'hb27;
      20'h00ebd: out <= 12'hf87;
      20'h00ebe: out <= 12'hf87;
      20'h00ebf: out <= 12'hf87;
      20'h00ec0: out <= 12'hf87;
      20'h00ec1: out <= 12'hf87;
      20'h00ec2: out <= 12'hf87;
      20'h00ec3: out <= 12'hee9;
      20'h00ec4: out <= 12'hb27;
      20'h00ec5: out <= 12'hf87;
      20'h00ec6: out <= 12'hf87;
      20'h00ec7: out <= 12'hf87;
      20'h00ec8: out <= 12'hf87;
      20'h00ec9: out <= 12'hf87;
      20'h00eca: out <= 12'hf87;
      20'h00ecb: out <= 12'hee9;
      20'h00ecc: out <= 12'h000;
      20'h00ecd: out <= 12'h000;
      20'h00ece: out <= 12'h000;
      20'h00ecf: out <= 12'h000;
      20'h00ed0: out <= 12'h000;
      20'h00ed1: out <= 12'h000;
      20'h00ed2: out <= 12'h000;
      20'h00ed3: out <= 12'h000;
      20'h00ed4: out <= 12'hb27;
      20'h00ed5: out <= 12'hf87;
      20'h00ed6: out <= 12'hf87;
      20'h00ed7: out <= 12'hf87;
      20'h00ed8: out <= 12'hf87;
      20'h00ed9: out <= 12'hf87;
      20'h00eda: out <= 12'hf87;
      20'h00edb: out <= 12'hee9;
      20'h00edc: out <= 12'hb27;
      20'h00edd: out <= 12'hf87;
      20'h00ede: out <= 12'hf87;
      20'h00edf: out <= 12'hf87;
      20'h00ee0: out <= 12'hf87;
      20'h00ee1: out <= 12'hf87;
      20'h00ee2: out <= 12'hf87;
      20'h00ee3: out <= 12'hee9;
      20'h00ee4: out <= 12'hb27;
      20'h00ee5: out <= 12'hf87;
      20'h00ee6: out <= 12'hf87;
      20'h00ee7: out <= 12'hf87;
      20'h00ee8: out <= 12'hf87;
      20'h00ee9: out <= 12'hf87;
      20'h00eea: out <= 12'hf87;
      20'h00eeb: out <= 12'hee9;
      20'h00eec: out <= 12'hb27;
      20'h00eed: out <= 12'hf87;
      20'h00eee: out <= 12'hf87;
      20'h00eef: out <= 12'hf87;
      20'h00ef0: out <= 12'hf87;
      20'h00ef1: out <= 12'hf87;
      20'h00ef2: out <= 12'hf87;
      20'h00ef3: out <= 12'hee9;
      20'h00ef4: out <= 12'h000;
      20'h00ef5: out <= 12'h000;
      20'h00ef6: out <= 12'h000;
      20'h00ef7: out <= 12'h000;
      20'h00ef8: out <= 12'h000;
      20'h00ef9: out <= 12'h000;
      20'h00efa: out <= 12'h000;
      20'h00efb: out <= 12'h000;
      20'h00efc: out <= 12'h000;
      20'h00efd: out <= 12'h000;
      20'h00efe: out <= 12'h000;
      20'h00eff: out <= 12'h000;
      20'h00f00: out <= 12'h000;
      20'h00f01: out <= 12'h000;
      20'h00f02: out <= 12'h000;
      20'h00f03: out <= 12'h000;
      20'h00f04: out <= 12'h000;
      20'h00f05: out <= 12'h000;
      20'h00f06: out <= 12'h000;
      20'h00f07: out <= 12'h000;
      20'h00f08: out <= 12'h000;
      20'h00f09: out <= 12'h000;
      20'h00f0a: out <= 12'h000;
      20'h00f0b: out <= 12'h000;
      20'h00f0c: out <= 12'h603;
      20'h00f0d: out <= 12'h603;
      20'h00f0e: out <= 12'h603;
      20'h00f0f: out <= 12'h603;
      20'h00f10: out <= 12'hee9;
      20'h00f11: out <= 12'hf87;
      20'h00f12: out <= 12'hee9;
      20'h00f13: out <= 12'hb27;
      20'h00f14: out <= 12'hb27;
      20'h00f15: out <= 12'hb27;
      20'h00f16: out <= 12'hf87;
      20'h00f17: out <= 12'hb27;
      20'h00f18: out <= 12'h000;
      20'h00f19: out <= 12'h000;
      20'h00f1a: out <= 12'h000;
      20'h00f1b: out <= 12'h000;
      20'h00f1c: out <= 12'h000;
      20'h00f1d: out <= 12'h000;
      20'h00f1e: out <= 12'h000;
      20'h00f1f: out <= 12'h000;
      20'h00f20: out <= 12'h000;
      20'h00f21: out <= 12'h000;
      20'h00f22: out <= 12'h000;
      20'h00f23: out <= 12'h000;
      20'h00f24: out <= 12'h000;
      20'h00f25: out <= 12'h000;
      20'h00f26: out <= 12'h000;
      20'h00f27: out <= 12'h000;
      20'h00f28: out <= 12'h000;
      20'h00f29: out <= 12'h000;
      20'h00f2a: out <= 12'h000;
      20'h00f2b: out <= 12'h000;
      20'h00f2c: out <= 12'h000;
      20'h00f2d: out <= 12'h000;
      20'h00f2e: out <= 12'h000;
      20'h00f2f: out <= 12'h000;
      20'h00f30: out <= 12'h000;
      20'h00f31: out <= 12'h000;
      20'h00f32: out <= 12'h000;
      20'h00f33: out <= 12'h000;
      20'h00f34: out <= 12'h000;
      20'h00f35: out <= 12'h000;
      20'h00f36: out <= 12'h000;
      20'h00f37: out <= 12'h000;
      20'h00f38: out <= 12'h000;
      20'h00f39: out <= 12'h000;
      20'h00f3a: out <= 12'h000;
      20'h00f3b: out <= 12'h000;
      20'h00f3c: out <= 12'h000;
      20'h00f3d: out <= 12'h000;
      20'h00f3e: out <= 12'h000;
      20'h00f3f: out <= 12'h000;
      20'h00f40: out <= 12'h000;
      20'h00f41: out <= 12'h000;
      20'h00f42: out <= 12'h000;
      20'h00f43: out <= 12'h000;
      20'h00f44: out <= 12'h000;
      20'h00f45: out <= 12'h000;
      20'h00f46: out <= 12'h000;
      20'h00f47: out <= 12'h000;
      20'h00f48: out <= 12'h000;
      20'h00f49: out <= 12'h000;
      20'h00f4a: out <= 12'h000;
      20'h00f4b: out <= 12'h000;
      20'h00f4c: out <= 12'h000;
      20'h00f4d: out <= 12'h000;
      20'h00f4e: out <= 12'h000;
      20'h00f4f: out <= 12'h000;
      20'h00f50: out <= 12'h222;
      20'h00f51: out <= 12'h6af;
      20'h00f52: out <= 12'h6af;
      20'h00f53: out <= 12'h6af;
      20'h00f54: out <= 12'h6af;
      20'h00f55: out <= 12'h6af;
      20'h00f56: out <= 12'h6af;
      20'h00f57: out <= 12'h6af;
      20'h00f58: out <= 12'h6af;
      20'h00f59: out <= 12'h6af;
      20'h00f5a: out <= 12'h6af;
      20'h00f5b: out <= 12'h6af;
      20'h00f5c: out <= 12'h6af;
      20'h00f5d: out <= 12'h222;
      20'h00f5e: out <= 12'h222;
      20'h00f5f: out <= 12'h222;
      20'h00f60: out <= 12'h000;
      20'h00f61: out <= 12'h6af;
      20'h00f62: out <= 12'h6af;
      20'h00f63: out <= 12'h6af;
      20'h00f64: out <= 12'h6af;
      20'h00f65: out <= 12'h6af;
      20'h00f66: out <= 12'h6af;
      20'h00f67: out <= 12'h6af;
      20'h00f68: out <= 12'h6af;
      20'h00f69: out <= 12'h6af;
      20'h00f6a: out <= 12'h6af;
      20'h00f6b: out <= 12'h6af;
      20'h00f6c: out <= 12'h6af;
      20'h00f6d: out <= 12'h000;
      20'h00f6e: out <= 12'h000;
      20'h00f6f: out <= 12'h000;
      20'h00f70: out <= 12'h222;
      20'h00f71: out <= 12'h6af;
      20'h00f72: out <= 12'hfff;
      20'h00f73: out <= 12'h6af;
      20'h00f74: out <= 12'h222;
      20'h00f75: out <= 12'h222;
      20'h00f76: out <= 12'h222;
      20'h00f77: out <= 12'h222;
      20'h00f78: out <= 12'h222;
      20'h00f79: out <= 12'h222;
      20'h00f7a: out <= 12'h222;
      20'h00f7b: out <= 12'h222;
      20'h00f7c: out <= 12'h222;
      20'h00f7d: out <= 12'h6af;
      20'h00f7e: out <= 12'hfff;
      20'h00f7f: out <= 12'h6af;
      20'h00f80: out <= 12'h000;
      20'h00f81: out <= 12'h6af;
      20'h00f82: out <= 12'h6af;
      20'h00f83: out <= 12'h6af;
      20'h00f84: out <= 12'h000;
      20'h00f85: out <= 12'h000;
      20'h00f86: out <= 12'h000;
      20'h00f87: out <= 12'h000;
      20'h00f88: out <= 12'h000;
      20'h00f89: out <= 12'h000;
      20'h00f8a: out <= 12'h000;
      20'h00f8b: out <= 12'h000;
      20'h00f8c: out <= 12'h000;
      20'h00f8d: out <= 12'h6af;
      20'h00f8e: out <= 12'h6af;
      20'h00f8f: out <= 12'h6af;
      20'h00f90: out <= 12'h222;
      20'h00f91: out <= 12'h222;
      20'h00f92: out <= 12'h222;
      20'h00f93: out <= 12'h6af;
      20'h00f94: out <= 12'h6af;
      20'h00f95: out <= 12'h6af;
      20'h00f96: out <= 12'h6af;
      20'h00f97: out <= 12'h6af;
      20'h00f98: out <= 12'h6af;
      20'h00f99: out <= 12'h6af;
      20'h00f9a: out <= 12'h6af;
      20'h00f9b: out <= 12'h6af;
      20'h00f9c: out <= 12'h6af;
      20'h00f9d: out <= 12'h6af;
      20'h00f9e: out <= 12'h6af;
      20'h00f9f: out <= 12'h222;
      20'h00fa0: out <= 12'h000;
      20'h00fa1: out <= 12'h000;
      20'h00fa2: out <= 12'h000;
      20'h00fa3: out <= 12'h6af;
      20'h00fa4: out <= 12'h6af;
      20'h00fa5: out <= 12'h6af;
      20'h00fa6: out <= 12'h6af;
      20'h00fa7: out <= 12'h6af;
      20'h00fa8: out <= 12'h6af;
      20'h00fa9: out <= 12'h6af;
      20'h00faa: out <= 12'h6af;
      20'h00fab: out <= 12'h6af;
      20'h00fac: out <= 12'h6af;
      20'h00fad: out <= 12'h6af;
      20'h00fae: out <= 12'h6af;
      20'h00faf: out <= 12'h000;
      20'h00fb0: out <= 12'h222;
      20'h00fb1: out <= 12'h222;
      20'h00fb2: out <= 12'h222;
      20'h00fb3: out <= 12'h222;
      20'h00fb4: out <= 12'h222;
      20'h00fb5: out <= 12'h222;
      20'h00fb6: out <= 12'h222;
      20'h00fb7: out <= 12'h16d;
      20'h00fb8: out <= 12'hfff;
      20'h00fb9: out <= 12'h16d;
      20'h00fba: out <= 12'h222;
      20'h00fbb: out <= 12'h222;
      20'h00fbc: out <= 12'h222;
      20'h00fbd: out <= 12'h222;
      20'h00fbe: out <= 12'h222;
      20'h00fbf: out <= 12'h222;
      20'h00fc0: out <= 12'h000;
      20'h00fc1: out <= 12'h000;
      20'h00fc2: out <= 12'h000;
      20'h00fc3: out <= 12'h000;
      20'h00fc4: out <= 12'h000;
      20'h00fc5: out <= 12'h000;
      20'h00fc6: out <= 12'h000;
      20'h00fc7: out <= 12'h16d;
      20'h00fc8: out <= 12'hfff;
      20'h00fc9: out <= 12'h16d;
      20'h00fca: out <= 12'h000;
      20'h00fcb: out <= 12'h000;
      20'h00fcc: out <= 12'h000;
      20'h00fcd: out <= 12'h000;
      20'h00fce: out <= 12'h000;
      20'h00fcf: out <= 12'h000;
      20'h00fd0: out <= 12'h603;
      20'h00fd1: out <= 12'h603;
      20'h00fd2: out <= 12'h603;
      20'h00fd3: out <= 12'h603;
      20'h00fd4: out <= 12'hb27;
      20'h00fd5: out <= 12'hf87;
      20'h00fd6: out <= 12'hf87;
      20'h00fd7: out <= 12'hf87;
      20'h00fd8: out <= 12'hf87;
      20'h00fd9: out <= 12'hf87;
      20'h00fda: out <= 12'hf87;
      20'h00fdb: out <= 12'hee9;
      20'h00fdc: out <= 12'hb27;
      20'h00fdd: out <= 12'hf87;
      20'h00fde: out <= 12'hf87;
      20'h00fdf: out <= 12'hf87;
      20'h00fe0: out <= 12'hf87;
      20'h00fe1: out <= 12'hf87;
      20'h00fe2: out <= 12'hf87;
      20'h00fe3: out <= 12'hee9;
      20'h00fe4: out <= 12'h000;
      20'h00fe5: out <= 12'h000;
      20'h00fe6: out <= 12'h000;
      20'h00fe7: out <= 12'h000;
      20'h00fe8: out <= 12'h000;
      20'h00fe9: out <= 12'h000;
      20'h00fea: out <= 12'h000;
      20'h00feb: out <= 12'h000;
      20'h00fec: out <= 12'hb27;
      20'h00fed: out <= 12'hf87;
      20'h00fee: out <= 12'hf87;
      20'h00fef: out <= 12'hf87;
      20'h00ff0: out <= 12'hf87;
      20'h00ff1: out <= 12'hf87;
      20'h00ff2: out <= 12'hf87;
      20'h00ff3: out <= 12'hee9;
      20'h00ff4: out <= 12'hb27;
      20'h00ff5: out <= 12'hf87;
      20'h00ff6: out <= 12'hf87;
      20'h00ff7: out <= 12'hf87;
      20'h00ff8: out <= 12'hf87;
      20'h00ff9: out <= 12'hf87;
      20'h00ffa: out <= 12'hf87;
      20'h00ffb: out <= 12'hee9;
      20'h00ffc: out <= 12'hb27;
      20'h00ffd: out <= 12'hf87;
      20'h00ffe: out <= 12'hf87;
      20'h00fff: out <= 12'hf87;
      20'h01000: out <= 12'hf87;
      20'h01001: out <= 12'hf87;
      20'h01002: out <= 12'hf87;
      20'h01003: out <= 12'hee9;
      20'h01004: out <= 12'hb27;
      20'h01005: out <= 12'hf87;
      20'h01006: out <= 12'hf87;
      20'h01007: out <= 12'hf87;
      20'h01008: out <= 12'hf87;
      20'h01009: out <= 12'hf87;
      20'h0100a: out <= 12'hf87;
      20'h0100b: out <= 12'hee9;
      20'h0100c: out <= 12'h000;
      20'h0100d: out <= 12'h000;
      20'h0100e: out <= 12'h000;
      20'h0100f: out <= 12'h000;
      20'h01010: out <= 12'h000;
      20'h01011: out <= 12'h000;
      20'h01012: out <= 12'h000;
      20'h01013: out <= 12'h000;
      20'h01014: out <= 12'h000;
      20'h01015: out <= 12'h000;
      20'h01016: out <= 12'h000;
      20'h01017: out <= 12'h000;
      20'h01018: out <= 12'h000;
      20'h01019: out <= 12'h000;
      20'h0101a: out <= 12'h000;
      20'h0101b: out <= 12'h000;
      20'h0101c: out <= 12'h000;
      20'h0101d: out <= 12'h000;
      20'h0101e: out <= 12'h000;
      20'h0101f: out <= 12'h000;
      20'h01020: out <= 12'h000;
      20'h01021: out <= 12'h000;
      20'h01022: out <= 12'h000;
      20'h01023: out <= 12'h000;
      20'h01024: out <= 12'h603;
      20'h01025: out <= 12'h603;
      20'h01026: out <= 12'h603;
      20'h01027: out <= 12'h603;
      20'h01028: out <= 12'hee9;
      20'h01029: out <= 12'hf87;
      20'h0102a: out <= 12'hf87;
      20'h0102b: out <= 12'hf87;
      20'h0102c: out <= 12'hf87;
      20'h0102d: out <= 12'hf87;
      20'h0102e: out <= 12'hf87;
      20'h0102f: out <= 12'hb27;
      20'h01030: out <= 12'h000;
      20'h01031: out <= 12'h000;
      20'h01032: out <= 12'h000;
      20'h01033: out <= 12'h000;
      20'h01034: out <= 12'h000;
      20'h01035: out <= 12'h000;
      20'h01036: out <= 12'h000;
      20'h01037: out <= 12'h000;
      20'h01038: out <= 12'h000;
      20'h01039: out <= 12'h000;
      20'h0103a: out <= 12'h000;
      20'h0103b: out <= 12'h000;
      20'h0103c: out <= 12'h000;
      20'h0103d: out <= 12'h000;
      20'h0103e: out <= 12'h000;
      20'h0103f: out <= 12'h000;
      20'h01040: out <= 12'h000;
      20'h01041: out <= 12'h000;
      20'h01042: out <= 12'h000;
      20'h01043: out <= 12'h000;
      20'h01044: out <= 12'h000;
      20'h01045: out <= 12'h000;
      20'h01046: out <= 12'h000;
      20'h01047: out <= 12'h000;
      20'h01048: out <= 12'h000;
      20'h01049: out <= 12'h000;
      20'h0104a: out <= 12'h000;
      20'h0104b: out <= 12'h000;
      20'h0104c: out <= 12'h000;
      20'h0104d: out <= 12'h000;
      20'h0104e: out <= 12'h000;
      20'h0104f: out <= 12'h000;
      20'h01050: out <= 12'h000;
      20'h01051: out <= 12'h000;
      20'h01052: out <= 12'h000;
      20'h01053: out <= 12'h000;
      20'h01054: out <= 12'h000;
      20'h01055: out <= 12'h000;
      20'h01056: out <= 12'h000;
      20'h01057: out <= 12'h000;
      20'h01058: out <= 12'h000;
      20'h01059: out <= 12'h000;
      20'h0105a: out <= 12'h000;
      20'h0105b: out <= 12'h000;
      20'h0105c: out <= 12'h000;
      20'h0105d: out <= 12'h000;
      20'h0105e: out <= 12'h000;
      20'h0105f: out <= 12'h000;
      20'h01060: out <= 12'h000;
      20'h01061: out <= 12'h000;
      20'h01062: out <= 12'h000;
      20'h01063: out <= 12'h000;
      20'h01064: out <= 12'h000;
      20'h01065: out <= 12'h000;
      20'h01066: out <= 12'h000;
      20'h01067: out <= 12'h000;
      20'h01068: out <= 12'h222;
      20'h01069: out <= 12'h222;
      20'h0106a: out <= 12'h222;
      20'h0106b: out <= 12'h222;
      20'h0106c: out <= 12'h222;
      20'h0106d: out <= 12'h222;
      20'h0106e: out <= 12'h222;
      20'h0106f: out <= 12'h222;
      20'h01070: out <= 12'h222;
      20'h01071: out <= 12'h222;
      20'h01072: out <= 12'h222;
      20'h01073: out <= 12'h222;
      20'h01074: out <= 12'h222;
      20'h01075: out <= 12'h222;
      20'h01076: out <= 12'h222;
      20'h01077: out <= 12'h222;
      20'h01078: out <= 12'h000;
      20'h01079: out <= 12'h000;
      20'h0107a: out <= 12'h000;
      20'h0107b: out <= 12'h000;
      20'h0107c: out <= 12'h000;
      20'h0107d: out <= 12'h000;
      20'h0107e: out <= 12'h000;
      20'h0107f: out <= 12'h000;
      20'h01080: out <= 12'h000;
      20'h01081: out <= 12'h000;
      20'h01082: out <= 12'h000;
      20'h01083: out <= 12'h000;
      20'h01084: out <= 12'h000;
      20'h01085: out <= 12'h000;
      20'h01086: out <= 12'h000;
      20'h01087: out <= 12'h000;
      20'h01088: out <= 12'h222;
      20'h01089: out <= 12'h222;
      20'h0108a: out <= 12'h222;
      20'h0108b: out <= 12'h222;
      20'h0108c: out <= 12'h222;
      20'h0108d: out <= 12'h222;
      20'h0108e: out <= 12'h222;
      20'h0108f: out <= 12'h222;
      20'h01090: out <= 12'h222;
      20'h01091: out <= 12'h222;
      20'h01092: out <= 12'h222;
      20'h01093: out <= 12'h222;
      20'h01094: out <= 12'h222;
      20'h01095: out <= 12'h222;
      20'h01096: out <= 12'h222;
      20'h01097: out <= 12'h222;
      20'h01098: out <= 12'h000;
      20'h01099: out <= 12'h000;
      20'h0109a: out <= 12'h000;
      20'h0109b: out <= 12'h000;
      20'h0109c: out <= 12'h000;
      20'h0109d: out <= 12'h000;
      20'h0109e: out <= 12'h000;
      20'h0109f: out <= 12'h000;
      20'h010a0: out <= 12'h000;
      20'h010a1: out <= 12'h000;
      20'h010a2: out <= 12'h000;
      20'h010a3: out <= 12'h000;
      20'h010a4: out <= 12'h000;
      20'h010a5: out <= 12'h000;
      20'h010a6: out <= 12'h000;
      20'h010a7: out <= 12'h000;
      20'h010a8: out <= 12'h222;
      20'h010a9: out <= 12'h222;
      20'h010aa: out <= 12'h222;
      20'h010ab: out <= 12'h222;
      20'h010ac: out <= 12'h222;
      20'h010ad: out <= 12'h222;
      20'h010ae: out <= 12'h222;
      20'h010af: out <= 12'h222;
      20'h010b0: out <= 12'h222;
      20'h010b1: out <= 12'h222;
      20'h010b2: out <= 12'h222;
      20'h010b3: out <= 12'h222;
      20'h010b4: out <= 12'h222;
      20'h010b5: out <= 12'h222;
      20'h010b6: out <= 12'h222;
      20'h010b7: out <= 12'h222;
      20'h010b8: out <= 12'h000;
      20'h010b9: out <= 12'h000;
      20'h010ba: out <= 12'h000;
      20'h010bb: out <= 12'h000;
      20'h010bc: out <= 12'h000;
      20'h010bd: out <= 12'h000;
      20'h010be: out <= 12'h000;
      20'h010bf: out <= 12'h000;
      20'h010c0: out <= 12'h000;
      20'h010c1: out <= 12'h000;
      20'h010c2: out <= 12'h000;
      20'h010c3: out <= 12'h000;
      20'h010c4: out <= 12'h000;
      20'h010c5: out <= 12'h000;
      20'h010c6: out <= 12'h000;
      20'h010c7: out <= 12'h000;
      20'h010c8: out <= 12'h222;
      20'h010c9: out <= 12'h222;
      20'h010ca: out <= 12'h222;
      20'h010cb: out <= 12'h222;
      20'h010cc: out <= 12'h222;
      20'h010cd: out <= 12'h222;
      20'h010ce: out <= 12'h222;
      20'h010cf: out <= 12'h6af;
      20'h010d0: out <= 12'hfff;
      20'h010d1: out <= 12'h6af;
      20'h010d2: out <= 12'h222;
      20'h010d3: out <= 12'h222;
      20'h010d4: out <= 12'h222;
      20'h010d5: out <= 12'h222;
      20'h010d6: out <= 12'h222;
      20'h010d7: out <= 12'h222;
      20'h010d8: out <= 12'h000;
      20'h010d9: out <= 12'h000;
      20'h010da: out <= 12'h000;
      20'h010db: out <= 12'h000;
      20'h010dc: out <= 12'h000;
      20'h010dd: out <= 12'h000;
      20'h010de: out <= 12'h000;
      20'h010df: out <= 12'h6af;
      20'h010e0: out <= 12'hfff;
      20'h010e1: out <= 12'h6af;
      20'h010e2: out <= 12'h000;
      20'h010e3: out <= 12'h000;
      20'h010e4: out <= 12'h000;
      20'h010e5: out <= 12'h000;
      20'h010e6: out <= 12'h000;
      20'h010e7: out <= 12'h000;
      20'h010e8: out <= 12'h603;
      20'h010e9: out <= 12'h603;
      20'h010ea: out <= 12'h603;
      20'h010eb: out <= 12'h603;
      20'h010ec: out <= 12'hb27;
      20'h010ed: out <= 12'hb27;
      20'h010ee: out <= 12'hb27;
      20'h010ef: out <= 12'hb27;
      20'h010f0: out <= 12'hb27;
      20'h010f1: out <= 12'hb27;
      20'h010f2: out <= 12'hb27;
      20'h010f3: out <= 12'hb27;
      20'h010f4: out <= 12'hb27;
      20'h010f5: out <= 12'hb27;
      20'h010f6: out <= 12'hb27;
      20'h010f7: out <= 12'hb27;
      20'h010f8: out <= 12'hb27;
      20'h010f9: out <= 12'hb27;
      20'h010fa: out <= 12'hb27;
      20'h010fb: out <= 12'hb27;
      20'h010fc: out <= 12'h000;
      20'h010fd: out <= 12'h000;
      20'h010fe: out <= 12'h000;
      20'h010ff: out <= 12'h000;
      20'h01100: out <= 12'h000;
      20'h01101: out <= 12'h000;
      20'h01102: out <= 12'h000;
      20'h01103: out <= 12'h000;
      20'h01104: out <= 12'hb27;
      20'h01105: out <= 12'hb27;
      20'h01106: out <= 12'hb27;
      20'h01107: out <= 12'hb27;
      20'h01108: out <= 12'hb27;
      20'h01109: out <= 12'hb27;
      20'h0110a: out <= 12'hb27;
      20'h0110b: out <= 12'hb27;
      20'h0110c: out <= 12'hb27;
      20'h0110d: out <= 12'hb27;
      20'h0110e: out <= 12'hb27;
      20'h0110f: out <= 12'hb27;
      20'h01110: out <= 12'hb27;
      20'h01111: out <= 12'hb27;
      20'h01112: out <= 12'hb27;
      20'h01113: out <= 12'hb27;
      20'h01114: out <= 12'hb27;
      20'h01115: out <= 12'hb27;
      20'h01116: out <= 12'hb27;
      20'h01117: out <= 12'hb27;
      20'h01118: out <= 12'hb27;
      20'h01119: out <= 12'hb27;
      20'h0111a: out <= 12'hb27;
      20'h0111b: out <= 12'hb27;
      20'h0111c: out <= 12'hb27;
      20'h0111d: out <= 12'hb27;
      20'h0111e: out <= 12'hb27;
      20'h0111f: out <= 12'hb27;
      20'h01120: out <= 12'hb27;
      20'h01121: out <= 12'hb27;
      20'h01122: out <= 12'hb27;
      20'h01123: out <= 12'hb27;
      20'h01124: out <= 12'h000;
      20'h01125: out <= 12'h000;
      20'h01126: out <= 12'h000;
      20'h01127: out <= 12'h000;
      20'h01128: out <= 12'h000;
      20'h01129: out <= 12'h000;
      20'h0112a: out <= 12'h000;
      20'h0112b: out <= 12'h000;
      20'h0112c: out <= 12'h000;
      20'h0112d: out <= 12'h000;
      20'h0112e: out <= 12'h000;
      20'h0112f: out <= 12'h000;
      20'h01130: out <= 12'h000;
      20'h01131: out <= 12'h000;
      20'h01132: out <= 12'h000;
      20'h01133: out <= 12'h000;
      20'h01134: out <= 12'h000;
      20'h01135: out <= 12'h000;
      20'h01136: out <= 12'h000;
      20'h01137: out <= 12'h000;
      20'h01138: out <= 12'h000;
      20'h01139: out <= 12'h000;
      20'h0113a: out <= 12'h000;
      20'h0113b: out <= 12'h000;
      20'h0113c: out <= 12'h603;
      20'h0113d: out <= 12'h603;
      20'h0113e: out <= 12'h603;
      20'h0113f: out <= 12'h603;
      20'h01140: out <= 12'hb27;
      20'h01141: out <= 12'hb27;
      20'h01142: out <= 12'hb27;
      20'h01143: out <= 12'hb27;
      20'h01144: out <= 12'hb27;
      20'h01145: out <= 12'hb27;
      20'h01146: out <= 12'hb27;
      20'h01147: out <= 12'hb27;
      20'h01148: out <= 12'h000;
      20'h01149: out <= 12'h000;
      20'h0114a: out <= 12'h000;
      20'h0114b: out <= 12'h000;
      20'h0114c: out <= 12'h000;
      20'h0114d: out <= 12'h000;
      20'h0114e: out <= 12'h000;
      20'h0114f: out <= 12'h000;
      20'h01150: out <= 12'h000;
      20'h01151: out <= 12'h000;
      20'h01152: out <= 12'h000;
      20'h01153: out <= 12'h000;
      20'h01154: out <= 12'h000;
      20'h01155: out <= 12'h000;
      20'h01156: out <= 12'h000;
      20'h01157: out <= 12'h000;
      20'h01158: out <= 12'h000;
      20'h01159: out <= 12'h000;
      20'h0115a: out <= 12'h000;
      20'h0115b: out <= 12'h000;
      20'h0115c: out <= 12'h000;
      20'h0115d: out <= 12'h000;
      20'h0115e: out <= 12'h000;
      20'h0115f: out <= 12'h000;
      20'h01160: out <= 12'h000;
      20'h01161: out <= 12'h000;
      20'h01162: out <= 12'h000;
      20'h01163: out <= 12'h000;
      20'h01164: out <= 12'h000;
      20'h01165: out <= 12'h000;
      20'h01166: out <= 12'h000;
      20'h01167: out <= 12'h000;
      20'h01168: out <= 12'h000;
      20'h01169: out <= 12'h000;
      20'h0116a: out <= 12'h000;
      20'h0116b: out <= 12'h000;
      20'h0116c: out <= 12'h000;
      20'h0116d: out <= 12'h000;
      20'h0116e: out <= 12'h000;
      20'h0116f: out <= 12'h000;
      20'h01170: out <= 12'h000;
      20'h01171: out <= 12'h000;
      20'h01172: out <= 12'h000;
      20'h01173: out <= 12'h000;
      20'h01174: out <= 12'h000;
      20'h01175: out <= 12'h000;
      20'h01176: out <= 12'h000;
      20'h01177: out <= 12'h000;
      20'h01178: out <= 12'h000;
      20'h01179: out <= 12'h000;
      20'h0117a: out <= 12'h000;
      20'h0117b: out <= 12'h000;
      20'h0117c: out <= 12'h000;
      20'h0117d: out <= 12'h000;
      20'h0117e: out <= 12'h000;
      20'h0117f: out <= 12'h000;
      20'h01180: out <= 12'h000;
      20'h01181: out <= 12'h6af;
      20'h01182: out <= 12'hfff;
      20'h01183: out <= 12'h6af;
      20'h01184: out <= 12'hfff;
      20'h01185: out <= 12'hfff;
      20'h01186: out <= 12'hfff;
      20'h01187: out <= 12'hfff;
      20'h01188: out <= 12'hfff;
      20'h01189: out <= 12'h6af;
      20'h0118a: out <= 12'h6af;
      20'h0118b: out <= 12'hfff;
      20'h0118c: out <= 12'h6af;
      20'h0118d: out <= 12'h000;
      20'h0118e: out <= 12'h000;
      20'h0118f: out <= 12'h000;
      20'h01190: out <= 12'h222;
      20'h01191: out <= 12'h6af;
      20'h01192: out <= 12'hfff;
      20'h01193: out <= 12'h6af;
      20'h01194: out <= 12'h16d;
      20'h01195: out <= 12'h16d;
      20'h01196: out <= 12'h16d;
      20'h01197: out <= 12'h16d;
      20'h01198: out <= 12'h16d;
      20'h01199: out <= 12'h6af;
      20'h0119a: out <= 12'h6af;
      20'h0119b: out <= 12'hfff;
      20'h0119c: out <= 12'h6af;
      20'h0119d: out <= 12'h222;
      20'h0119e: out <= 12'h222;
      20'h0119f: out <= 12'h222;
      20'h011a0: out <= 12'h000;
      20'h011a1: out <= 12'h000;
      20'h011a2: out <= 12'h000;
      20'h011a3: out <= 12'h000;
      20'h011a4: out <= 12'h000;
      20'h011a5: out <= 12'h000;
      20'h011a6: out <= 12'h000;
      20'h011a7: out <= 12'h6af;
      20'h011a8: out <= 12'hfff;
      20'h011a9: out <= 12'h6af;
      20'h011aa: out <= 12'h000;
      20'h011ab: out <= 12'h000;
      20'h011ac: out <= 12'h000;
      20'h011ad: out <= 12'h000;
      20'h011ae: out <= 12'h000;
      20'h011af: out <= 12'h000;
      20'h011b0: out <= 12'h222;
      20'h011b1: out <= 12'h222;
      20'h011b2: out <= 12'h222;
      20'h011b3: out <= 12'h222;
      20'h011b4: out <= 12'h222;
      20'h011b5: out <= 12'h222;
      20'h011b6: out <= 12'h222;
      20'h011b7: out <= 12'h6af;
      20'h011b8: out <= 12'hfff;
      20'h011b9: out <= 12'h6af;
      20'h011ba: out <= 12'h222;
      20'h011bb: out <= 12'h222;
      20'h011bc: out <= 12'h222;
      20'h011bd: out <= 12'h222;
      20'h011be: out <= 12'h222;
      20'h011bf: out <= 12'h222;
      20'h011c0: out <= 12'h000;
      20'h011c1: out <= 12'h000;
      20'h011c2: out <= 12'h000;
      20'h011c3: out <= 12'h6af;
      20'h011c4: out <= 12'hfff;
      20'h011c5: out <= 12'h6af;
      20'h011c6: out <= 12'h6af;
      20'h011c7: out <= 12'hfff;
      20'h011c8: out <= 12'hfff;
      20'h011c9: out <= 12'hfff;
      20'h011ca: out <= 12'hfff;
      20'h011cb: out <= 12'hfff;
      20'h011cc: out <= 12'h6af;
      20'h011cd: out <= 12'hfff;
      20'h011ce: out <= 12'h6af;
      20'h011cf: out <= 12'h000;
      20'h011d0: out <= 12'h222;
      20'h011d1: out <= 12'h222;
      20'h011d2: out <= 12'h222;
      20'h011d3: out <= 12'h6af;
      20'h011d4: out <= 12'hfff;
      20'h011d5: out <= 12'h6af;
      20'h011d6: out <= 12'h6af;
      20'h011d7: out <= 12'h16d;
      20'h011d8: out <= 12'h16d;
      20'h011d9: out <= 12'h16d;
      20'h011da: out <= 12'h16d;
      20'h011db: out <= 12'h16d;
      20'h011dc: out <= 12'h6af;
      20'h011dd: out <= 12'hfff;
      20'h011de: out <= 12'h6af;
      20'h011df: out <= 12'h222;
      20'h011e0: out <= 12'h000;
      20'h011e1: out <= 12'h000;
      20'h011e2: out <= 12'h000;
      20'h011e3: out <= 12'h000;
      20'h011e4: out <= 12'h000;
      20'h011e5: out <= 12'h000;
      20'h011e6: out <= 12'hfff;
      20'h011e7: out <= 12'hfff;
      20'h011e8: out <= 12'hfff;
      20'h011e9: out <= 12'hfff;
      20'h011ea: out <= 12'hfff;
      20'h011eb: out <= 12'h000;
      20'h011ec: out <= 12'h000;
      20'h011ed: out <= 12'h000;
      20'h011ee: out <= 12'h000;
      20'h011ef: out <= 12'h000;
      20'h011f0: out <= 12'h222;
      20'h011f1: out <= 12'h222;
      20'h011f2: out <= 12'h222;
      20'h011f3: out <= 12'h222;
      20'h011f4: out <= 12'h222;
      20'h011f5: out <= 12'h222;
      20'h011f6: out <= 12'h16d;
      20'h011f7: out <= 12'h16d;
      20'h011f8: out <= 12'h16d;
      20'h011f9: out <= 12'h16d;
      20'h011fa: out <= 12'h16d;
      20'h011fb: out <= 12'h222;
      20'h011fc: out <= 12'h222;
      20'h011fd: out <= 12'h222;
      20'h011fe: out <= 12'h222;
      20'h011ff: out <= 12'h222;
      20'h01200: out <= 12'h603;
      20'h01201: out <= 12'h603;
      20'h01202: out <= 12'h603;
      20'h01203: out <= 12'h603;
      20'h01204: out <= 12'hfff;
      20'h01205: out <= 12'hfff;
      20'h01206: out <= 12'hfff;
      20'h01207: out <= 12'hfff;
      20'h01208: out <= 12'hfff;
      20'h01209: out <= 12'hfff;
      20'h0120a: out <= 12'hfff;
      20'h0120b: out <= 12'h666;
      20'h0120c: out <= 12'hfff;
      20'h0120d: out <= 12'hfff;
      20'h0120e: out <= 12'hfff;
      20'h0120f: out <= 12'hfff;
      20'h01210: out <= 12'hfff;
      20'h01211: out <= 12'hfff;
      20'h01212: out <= 12'hfff;
      20'h01213: out <= 12'h666;
      20'h01214: out <= 12'h000;
      20'h01215: out <= 12'h000;
      20'h01216: out <= 12'h000;
      20'h01217: out <= 12'h000;
      20'h01218: out <= 12'h000;
      20'h01219: out <= 12'h000;
      20'h0121a: out <= 12'h000;
      20'h0121b: out <= 12'h000;
      20'h0121c: out <= 12'hfff;
      20'h0121d: out <= 12'hfff;
      20'h0121e: out <= 12'hfff;
      20'h0121f: out <= 12'hfff;
      20'h01220: out <= 12'hfff;
      20'h01221: out <= 12'hfff;
      20'h01222: out <= 12'hfff;
      20'h01223: out <= 12'h666;
      20'h01224: out <= 12'h000;
      20'h01225: out <= 12'h000;
      20'h01226: out <= 12'h000;
      20'h01227: out <= 12'h000;
      20'h01228: out <= 12'h000;
      20'h01229: out <= 12'h000;
      20'h0122a: out <= 12'h000;
      20'h0122b: out <= 12'h000;
      20'h0122c: out <= 12'h000;
      20'h0122d: out <= 12'h000;
      20'h0122e: out <= 12'h000;
      20'h0122f: out <= 12'h000;
      20'h01230: out <= 12'h000;
      20'h01231: out <= 12'h000;
      20'h01232: out <= 12'h000;
      20'h01233: out <= 12'h000;
      20'h01234: out <= 12'hfff;
      20'h01235: out <= 12'hfff;
      20'h01236: out <= 12'hfff;
      20'h01237: out <= 12'hfff;
      20'h01238: out <= 12'hfff;
      20'h01239: out <= 12'hfff;
      20'h0123a: out <= 12'hfff;
      20'h0123b: out <= 12'h666;
      20'h0123c: out <= 12'h000;
      20'h0123d: out <= 12'h000;
      20'h0123e: out <= 12'h000;
      20'h0123f: out <= 12'h000;
      20'h01240: out <= 12'h000;
      20'h01241: out <= 12'h000;
      20'h01242: out <= 12'h000;
      20'h01243: out <= 12'h000;
      20'h01244: out <= 12'hfff;
      20'h01245: out <= 12'hfff;
      20'h01246: out <= 12'hfff;
      20'h01247: out <= 12'hfff;
      20'h01248: out <= 12'hfff;
      20'h01249: out <= 12'hfff;
      20'h0124a: out <= 12'hfff;
      20'h0124b: out <= 12'h666;
      20'h0124c: out <= 12'hfff;
      20'h0124d: out <= 12'hfff;
      20'h0124e: out <= 12'hfff;
      20'h0124f: out <= 12'hfff;
      20'h01250: out <= 12'hfff;
      20'h01251: out <= 12'hfff;
      20'h01252: out <= 12'hfff;
      20'h01253: out <= 12'h666;
      20'h01254: out <= 12'h603;
      20'h01255: out <= 12'h603;
      20'h01256: out <= 12'h603;
      20'h01257: out <= 12'h603;
      20'h01258: out <= 12'hee9;
      20'h01259: out <= 12'hee9;
      20'h0125a: out <= 12'hee9;
      20'h0125b: out <= 12'hee9;
      20'h0125c: out <= 12'hee9;
      20'h0125d: out <= 12'hee9;
      20'h0125e: out <= 12'hee9;
      20'h0125f: out <= 12'hb27;
      20'h01260: out <= 12'h000;
      20'h01261: out <= 12'h000;
      20'h01262: out <= 12'h000;
      20'h01263: out <= 12'h000;
      20'h01264: out <= 12'h000;
      20'h01265: out <= 12'h000;
      20'h01266: out <= 12'h000;
      20'h01267: out <= 12'h000;
      20'h01268: out <= 12'h000;
      20'h01269: out <= 12'hee9;
      20'h0126a: out <= 12'hee9;
      20'h0126b: out <= 12'hee9;
      20'h0126c: out <= 12'hee9;
      20'h0126d: out <= 12'h000;
      20'h0126e: out <= 12'h000;
      20'h0126f: out <= 12'hee9;
      20'h01270: out <= 12'hee9;
      20'h01271: out <= 12'hee9;
      20'h01272: out <= 12'hee9;
      20'h01273: out <= 12'hee9;
      20'h01274: out <= 12'hee9;
      20'h01275: out <= 12'h000;
      20'h01276: out <= 12'h000;
      20'h01277: out <= 12'hee9;
      20'h01278: out <= 12'hee9;
      20'h01279: out <= 12'hee9;
      20'h0127a: out <= 12'hee9;
      20'h0127b: out <= 12'h000;
      20'h0127c: out <= 12'h000;
      20'h0127d: out <= 12'h000;
      20'h0127e: out <= 12'hee9;
      20'h0127f: out <= 12'hee9;
      20'h01280: out <= 12'hee9;
      20'h01281: out <= 12'hee9;
      20'h01282: out <= 12'h000;
      20'h01283: out <= 12'h000;
      20'h01284: out <= 12'hee9;
      20'h01285: out <= 12'hee9;
      20'h01286: out <= 12'hee9;
      20'h01287: out <= 12'hee9;
      20'h01288: out <= 12'hee9;
      20'h01289: out <= 12'h000;
      20'h0128a: out <= 12'h000;
      20'h0128b: out <= 12'h000;
      20'h0128c: out <= 12'h000;
      20'h0128d: out <= 12'h000;
      20'h0128e: out <= 12'h000;
      20'h0128f: out <= 12'h000;
      20'h01290: out <= 12'h000;
      20'h01291: out <= 12'h000;
      20'h01292: out <= 12'h000;
      20'h01293: out <= 12'h000;
      20'h01294: out <= 12'h000;
      20'h01295: out <= 12'h000;
      20'h01296: out <= 12'h000;
      20'h01297: out <= 12'h000;
      20'h01298: out <= 12'h000;
      20'h01299: out <= 12'h16d;
      20'h0129a: out <= 12'hfff;
      20'h0129b: out <= 12'hfff;
      20'h0129c: out <= 12'h6af;
      20'h0129d: out <= 12'h6af;
      20'h0129e: out <= 12'h6af;
      20'h0129f: out <= 12'h6af;
      20'h012a0: out <= 12'h6af;
      20'h012a1: out <= 12'hfff;
      20'h012a2: out <= 12'h16d;
      20'h012a3: out <= 12'hfff;
      20'h012a4: out <= 12'h16d;
      20'h012a5: out <= 12'h000;
      20'h012a6: out <= 12'h000;
      20'h012a7: out <= 12'h000;
      20'h012a8: out <= 12'h222;
      20'h012a9: out <= 12'h16d;
      20'h012aa: out <= 12'hfff;
      20'h012ab: out <= 12'h16d;
      20'h012ac: out <= 12'h6af;
      20'h012ad: out <= 12'h6af;
      20'h012ae: out <= 12'h6af;
      20'h012af: out <= 12'h6af;
      20'h012b0: out <= 12'h6af;
      20'h012b1: out <= 12'h16d;
      20'h012b2: out <= 12'h16d;
      20'h012b3: out <= 12'hfff;
      20'h012b4: out <= 12'h16d;
      20'h012b5: out <= 12'h222;
      20'h012b6: out <= 12'h222;
      20'h012b7: out <= 12'h222;
      20'h012b8: out <= 12'h000;
      20'h012b9: out <= 12'h000;
      20'h012ba: out <= 12'h000;
      20'h012bb: out <= 12'h000;
      20'h012bc: out <= 12'h000;
      20'h012bd: out <= 12'h000;
      20'h012be: out <= 12'h000;
      20'h012bf: out <= 12'h16d;
      20'h012c0: out <= 12'hfff;
      20'h012c1: out <= 12'h16d;
      20'h012c2: out <= 12'h000;
      20'h012c3: out <= 12'h000;
      20'h012c4: out <= 12'h000;
      20'h012c5: out <= 12'h000;
      20'h012c6: out <= 12'h000;
      20'h012c7: out <= 12'h000;
      20'h012c8: out <= 12'h222;
      20'h012c9: out <= 12'h222;
      20'h012ca: out <= 12'h222;
      20'h012cb: out <= 12'h222;
      20'h012cc: out <= 12'h222;
      20'h012cd: out <= 12'h222;
      20'h012ce: out <= 12'h222;
      20'h012cf: out <= 12'h16d;
      20'h012d0: out <= 12'hfff;
      20'h012d1: out <= 12'h16d;
      20'h012d2: out <= 12'h222;
      20'h012d3: out <= 12'h222;
      20'h012d4: out <= 12'h222;
      20'h012d5: out <= 12'h222;
      20'h012d6: out <= 12'h222;
      20'h012d7: out <= 12'h222;
      20'h012d8: out <= 12'h000;
      20'h012d9: out <= 12'h000;
      20'h012da: out <= 12'h000;
      20'h012db: out <= 12'h16d;
      20'h012dc: out <= 12'hfff;
      20'h012dd: out <= 12'h16d;
      20'h012de: out <= 12'hfff;
      20'h012df: out <= 12'h6af;
      20'h012e0: out <= 12'h6af;
      20'h012e1: out <= 12'h6af;
      20'h012e2: out <= 12'h6af;
      20'h012e3: out <= 12'h6af;
      20'h012e4: out <= 12'hfff;
      20'h012e5: out <= 12'hfff;
      20'h012e6: out <= 12'h16d;
      20'h012e7: out <= 12'h000;
      20'h012e8: out <= 12'h222;
      20'h012e9: out <= 12'h222;
      20'h012ea: out <= 12'h222;
      20'h012eb: out <= 12'h16d;
      20'h012ec: out <= 12'hfff;
      20'h012ed: out <= 12'h16d;
      20'h012ee: out <= 12'h16d;
      20'h012ef: out <= 12'h6af;
      20'h012f0: out <= 12'h6af;
      20'h012f1: out <= 12'h6af;
      20'h012f2: out <= 12'h6af;
      20'h012f3: out <= 12'h6af;
      20'h012f4: out <= 12'h16d;
      20'h012f5: out <= 12'hfff;
      20'h012f6: out <= 12'h16d;
      20'h012f7: out <= 12'h222;
      20'h012f8: out <= 12'h000;
      20'h012f9: out <= 12'h6af;
      20'h012fa: out <= 12'h16d;
      20'h012fb: out <= 12'h6af;
      20'h012fc: out <= 12'hfff;
      20'h012fd: out <= 12'hfff;
      20'h012fe: out <= 12'h6af;
      20'h012ff: out <= 12'h6af;
      20'h01300: out <= 12'h6af;
      20'h01301: out <= 12'h6af;
      20'h01302: out <= 12'h6af;
      20'h01303: out <= 12'hfff;
      20'h01304: out <= 12'hfff;
      20'h01305: out <= 12'h6af;
      20'h01306: out <= 12'h16d;
      20'h01307: out <= 12'h6af;
      20'h01308: out <= 12'h222;
      20'h01309: out <= 12'h6af;
      20'h0130a: out <= 12'h16d;
      20'h0130b: out <= 12'h6af;
      20'h0130c: out <= 12'h16d;
      20'h0130d: out <= 12'h16d;
      20'h0130e: out <= 12'h6af;
      20'h0130f: out <= 12'h6af;
      20'h01310: out <= 12'h6af;
      20'h01311: out <= 12'h6af;
      20'h01312: out <= 12'h6af;
      20'h01313: out <= 12'h16d;
      20'h01314: out <= 12'h16d;
      20'h01315: out <= 12'h6af;
      20'h01316: out <= 12'h16d;
      20'h01317: out <= 12'h6af;
      20'h01318: out <= 12'h603;
      20'h01319: out <= 12'h603;
      20'h0131a: out <= 12'h603;
      20'h0131b: out <= 12'h603;
      20'h0131c: out <= 12'hfff;
      20'h0131d: out <= 12'hbbb;
      20'h0131e: out <= 12'hbbb;
      20'h0131f: out <= 12'hbbb;
      20'h01320: out <= 12'hbbb;
      20'h01321: out <= 12'hbbb;
      20'h01322: out <= 12'h666;
      20'h01323: out <= 12'h666;
      20'h01324: out <= 12'hfff;
      20'h01325: out <= 12'hbbb;
      20'h01326: out <= 12'hbbb;
      20'h01327: out <= 12'hbbb;
      20'h01328: out <= 12'hbbb;
      20'h01329: out <= 12'hbbb;
      20'h0132a: out <= 12'h666;
      20'h0132b: out <= 12'h666;
      20'h0132c: out <= 12'h000;
      20'h0132d: out <= 12'h000;
      20'h0132e: out <= 12'h000;
      20'h0132f: out <= 12'h000;
      20'h01330: out <= 12'h000;
      20'h01331: out <= 12'h000;
      20'h01332: out <= 12'h000;
      20'h01333: out <= 12'h000;
      20'h01334: out <= 12'hfff;
      20'h01335: out <= 12'hbbb;
      20'h01336: out <= 12'hbbb;
      20'h01337: out <= 12'hbbb;
      20'h01338: out <= 12'hbbb;
      20'h01339: out <= 12'hbbb;
      20'h0133a: out <= 12'h666;
      20'h0133b: out <= 12'h666;
      20'h0133c: out <= 12'h000;
      20'h0133d: out <= 12'h000;
      20'h0133e: out <= 12'h000;
      20'h0133f: out <= 12'h000;
      20'h01340: out <= 12'h000;
      20'h01341: out <= 12'h000;
      20'h01342: out <= 12'h000;
      20'h01343: out <= 12'h000;
      20'h01344: out <= 12'h000;
      20'h01345: out <= 12'h000;
      20'h01346: out <= 12'h000;
      20'h01347: out <= 12'h000;
      20'h01348: out <= 12'h000;
      20'h01349: out <= 12'h000;
      20'h0134a: out <= 12'h000;
      20'h0134b: out <= 12'h000;
      20'h0134c: out <= 12'hfff;
      20'h0134d: out <= 12'hbbb;
      20'h0134e: out <= 12'hbbb;
      20'h0134f: out <= 12'hbbb;
      20'h01350: out <= 12'hbbb;
      20'h01351: out <= 12'hbbb;
      20'h01352: out <= 12'h666;
      20'h01353: out <= 12'h666;
      20'h01354: out <= 12'h000;
      20'h01355: out <= 12'h000;
      20'h01356: out <= 12'h000;
      20'h01357: out <= 12'h000;
      20'h01358: out <= 12'h000;
      20'h01359: out <= 12'h000;
      20'h0135a: out <= 12'h000;
      20'h0135b: out <= 12'h000;
      20'h0135c: out <= 12'hfff;
      20'h0135d: out <= 12'hbbb;
      20'h0135e: out <= 12'hbbb;
      20'h0135f: out <= 12'hbbb;
      20'h01360: out <= 12'hbbb;
      20'h01361: out <= 12'hbbb;
      20'h01362: out <= 12'h666;
      20'h01363: out <= 12'h666;
      20'h01364: out <= 12'hfff;
      20'h01365: out <= 12'hbbb;
      20'h01366: out <= 12'hbbb;
      20'h01367: out <= 12'hbbb;
      20'h01368: out <= 12'hbbb;
      20'h01369: out <= 12'hbbb;
      20'h0136a: out <= 12'h666;
      20'h0136b: out <= 12'h666;
      20'h0136c: out <= 12'h603;
      20'h0136d: out <= 12'h603;
      20'h0136e: out <= 12'h603;
      20'h0136f: out <= 12'h603;
      20'h01370: out <= 12'hee9;
      20'h01371: out <= 12'hf87;
      20'h01372: out <= 12'hf87;
      20'h01373: out <= 12'hf87;
      20'h01374: out <= 12'hf87;
      20'h01375: out <= 12'hf87;
      20'h01376: out <= 12'hf87;
      20'h01377: out <= 12'hb27;
      20'h01378: out <= 12'h000;
      20'h01379: out <= 12'h000;
      20'h0137a: out <= 12'h000;
      20'h0137b: out <= 12'h000;
      20'h0137c: out <= 12'h000;
      20'h0137d: out <= 12'h000;
      20'h0137e: out <= 12'h000;
      20'h0137f: out <= 12'h000;
      20'h01380: out <= 12'hee9;
      20'h01381: out <= 12'hee9;
      20'h01382: out <= 12'h000;
      20'h01383: out <= 12'h000;
      20'h01384: out <= 12'hee9;
      20'h01385: out <= 12'hee9;
      20'h01386: out <= 12'h000;
      20'h01387: out <= 12'h000;
      20'h01388: out <= 12'h000;
      20'h01389: out <= 12'hee9;
      20'h0138a: out <= 12'hee9;
      20'h0138b: out <= 12'h000;
      20'h0138c: out <= 12'h000;
      20'h0138d: out <= 12'h000;
      20'h0138e: out <= 12'hee9;
      20'h0138f: out <= 12'hee9;
      20'h01390: out <= 12'hee9;
      20'h01391: out <= 12'hee9;
      20'h01392: out <= 12'hee9;
      20'h01393: out <= 12'hee9;
      20'h01394: out <= 12'h000;
      20'h01395: out <= 12'hee9;
      20'h01396: out <= 12'hee9;
      20'h01397: out <= 12'h000;
      20'h01398: out <= 12'h000;
      20'h01399: out <= 12'hee9;
      20'h0139a: out <= 12'hee9;
      20'h0139b: out <= 12'h000;
      20'h0139c: out <= 12'hee9;
      20'h0139d: out <= 12'hee9;
      20'h0139e: out <= 12'h000;
      20'h0139f: out <= 12'h000;
      20'h013a0: out <= 12'h000;
      20'h013a1: out <= 12'h000;
      20'h013a2: out <= 12'h000;
      20'h013a3: out <= 12'h000;
      20'h013a4: out <= 12'h000;
      20'h013a5: out <= 12'h000;
      20'h013a6: out <= 12'h000;
      20'h013a7: out <= 12'h000;
      20'h013a8: out <= 12'h000;
      20'h013a9: out <= 12'h000;
      20'h013aa: out <= 12'h000;
      20'h013ab: out <= 12'h000;
      20'h013ac: out <= 12'h000;
      20'h013ad: out <= 12'h000;
      20'h013ae: out <= 12'h000;
      20'h013af: out <= 12'h000;
      20'h013b0: out <= 12'h000;
      20'h013b1: out <= 12'h6af;
      20'h013b2: out <= 12'hfff;
      20'h013b3: out <= 12'h6af;
      20'h013b4: out <= 12'h16d;
      20'h013b5: out <= 12'h16d;
      20'h013b6: out <= 12'h16d;
      20'h013b7: out <= 12'h16d;
      20'h013b8: out <= 12'h16d;
      20'h013b9: out <= 12'h6af;
      20'h013ba: out <= 12'hfff;
      20'h013bb: out <= 12'hfff;
      20'h013bc: out <= 12'h6af;
      20'h013bd: out <= 12'h000;
      20'h013be: out <= 12'h000;
      20'h013bf: out <= 12'h000;
      20'h013c0: out <= 12'h222;
      20'h013c1: out <= 12'h6af;
      20'h013c2: out <= 12'hfff;
      20'h013c3: out <= 12'h6af;
      20'h013c4: out <= 12'hfff;
      20'h013c5: out <= 12'hfff;
      20'h013c6: out <= 12'hfff;
      20'h013c7: out <= 12'hfff;
      20'h013c8: out <= 12'hfff;
      20'h013c9: out <= 12'h6af;
      20'h013ca: out <= 12'h16d;
      20'h013cb: out <= 12'hfff;
      20'h013cc: out <= 12'h6af;
      20'h013cd: out <= 12'h222;
      20'h013ce: out <= 12'h222;
      20'h013cf: out <= 12'h222;
      20'h013d0: out <= 12'h000;
      20'h013d1: out <= 12'h000;
      20'h013d2: out <= 12'h000;
      20'h013d3: out <= 12'h000;
      20'h013d4: out <= 12'h000;
      20'h013d5: out <= 12'h000;
      20'h013d6: out <= 12'h000;
      20'h013d7: out <= 12'h16d;
      20'h013d8: out <= 12'hfff;
      20'h013d9: out <= 12'h16d;
      20'h013da: out <= 12'h000;
      20'h013db: out <= 12'h000;
      20'h013dc: out <= 12'h000;
      20'h013dd: out <= 12'h000;
      20'h013de: out <= 12'h000;
      20'h013df: out <= 12'h000;
      20'h013e0: out <= 12'h222;
      20'h013e1: out <= 12'h222;
      20'h013e2: out <= 12'h222;
      20'h013e3: out <= 12'h222;
      20'h013e4: out <= 12'h222;
      20'h013e5: out <= 12'h222;
      20'h013e6: out <= 12'h222;
      20'h013e7: out <= 12'h16d;
      20'h013e8: out <= 12'hfff;
      20'h013e9: out <= 12'h16d;
      20'h013ea: out <= 12'h222;
      20'h013eb: out <= 12'h222;
      20'h013ec: out <= 12'h222;
      20'h013ed: out <= 12'h222;
      20'h013ee: out <= 12'h222;
      20'h013ef: out <= 12'h222;
      20'h013f0: out <= 12'h000;
      20'h013f1: out <= 12'h000;
      20'h013f2: out <= 12'h000;
      20'h013f3: out <= 12'h6af;
      20'h013f4: out <= 12'hfff;
      20'h013f5: out <= 12'hfff;
      20'h013f6: out <= 12'h6af;
      20'h013f7: out <= 12'h16d;
      20'h013f8: out <= 12'h16d;
      20'h013f9: out <= 12'h16d;
      20'h013fa: out <= 12'h16d;
      20'h013fb: out <= 12'h16d;
      20'h013fc: out <= 12'h6af;
      20'h013fd: out <= 12'hfff;
      20'h013fe: out <= 12'h6af;
      20'h013ff: out <= 12'h000;
      20'h01400: out <= 12'h222;
      20'h01401: out <= 12'h222;
      20'h01402: out <= 12'h222;
      20'h01403: out <= 12'h6af;
      20'h01404: out <= 12'hfff;
      20'h01405: out <= 12'h16d;
      20'h01406: out <= 12'h6af;
      20'h01407: out <= 12'hfff;
      20'h01408: out <= 12'hfff;
      20'h01409: out <= 12'hfff;
      20'h0140a: out <= 12'hfff;
      20'h0140b: out <= 12'hfff;
      20'h0140c: out <= 12'h6af;
      20'h0140d: out <= 12'hfff;
      20'h0140e: out <= 12'h6af;
      20'h0140f: out <= 12'h222;
      20'h01410: out <= 12'h000;
      20'h01411: out <= 12'hfff;
      20'h01412: out <= 12'hfff;
      20'h01413: out <= 12'hfff;
      20'h01414: out <= 12'h6af;
      20'h01415: out <= 12'h6af;
      20'h01416: out <= 12'h16d;
      20'h01417: out <= 12'h16d;
      20'h01418: out <= 12'h16d;
      20'h01419: out <= 12'h16d;
      20'h0141a: out <= 12'h16d;
      20'h0141b: out <= 12'h6af;
      20'h0141c: out <= 12'h6af;
      20'h0141d: out <= 12'hfff;
      20'h0141e: out <= 12'hfff;
      20'h0141f: out <= 12'hfff;
      20'h01420: out <= 12'h222;
      20'h01421: out <= 12'hfff;
      20'h01422: out <= 12'hfff;
      20'h01423: out <= 12'hfff;
      20'h01424: out <= 12'h6af;
      20'h01425: out <= 12'h6af;
      20'h01426: out <= 12'hfff;
      20'h01427: out <= 12'hfff;
      20'h01428: out <= 12'hfff;
      20'h01429: out <= 12'hfff;
      20'h0142a: out <= 12'hfff;
      20'h0142b: out <= 12'h6af;
      20'h0142c: out <= 12'h6af;
      20'h0142d: out <= 12'hfff;
      20'h0142e: out <= 12'hfff;
      20'h0142f: out <= 12'hfff;
      20'h01430: out <= 12'h603;
      20'h01431: out <= 12'h603;
      20'h01432: out <= 12'h603;
      20'h01433: out <= 12'h603;
      20'h01434: out <= 12'hfff;
      20'h01435: out <= 12'hbbb;
      20'h01436: out <= 12'h666;
      20'h01437: out <= 12'h666;
      20'h01438: out <= 12'h666;
      20'h01439: out <= 12'hbbb;
      20'h0143a: out <= 12'h666;
      20'h0143b: out <= 12'h666;
      20'h0143c: out <= 12'hfff;
      20'h0143d: out <= 12'hbbb;
      20'h0143e: out <= 12'h666;
      20'h0143f: out <= 12'h666;
      20'h01440: out <= 12'h666;
      20'h01441: out <= 12'hbbb;
      20'h01442: out <= 12'h666;
      20'h01443: out <= 12'h666;
      20'h01444: out <= 12'h000;
      20'h01445: out <= 12'h000;
      20'h01446: out <= 12'h000;
      20'h01447: out <= 12'h000;
      20'h01448: out <= 12'h000;
      20'h01449: out <= 12'h000;
      20'h0144a: out <= 12'h000;
      20'h0144b: out <= 12'h000;
      20'h0144c: out <= 12'hfff;
      20'h0144d: out <= 12'hbbb;
      20'h0144e: out <= 12'h666;
      20'h0144f: out <= 12'h666;
      20'h01450: out <= 12'h666;
      20'h01451: out <= 12'hbbb;
      20'h01452: out <= 12'h666;
      20'h01453: out <= 12'h666;
      20'h01454: out <= 12'h000;
      20'h01455: out <= 12'h000;
      20'h01456: out <= 12'h000;
      20'h01457: out <= 12'h000;
      20'h01458: out <= 12'h000;
      20'h01459: out <= 12'h000;
      20'h0145a: out <= 12'h000;
      20'h0145b: out <= 12'h000;
      20'h0145c: out <= 12'h000;
      20'h0145d: out <= 12'h000;
      20'h0145e: out <= 12'h000;
      20'h0145f: out <= 12'h000;
      20'h01460: out <= 12'h000;
      20'h01461: out <= 12'h000;
      20'h01462: out <= 12'h000;
      20'h01463: out <= 12'h000;
      20'h01464: out <= 12'hfff;
      20'h01465: out <= 12'hbbb;
      20'h01466: out <= 12'h666;
      20'h01467: out <= 12'h666;
      20'h01468: out <= 12'h666;
      20'h01469: out <= 12'hbbb;
      20'h0146a: out <= 12'h666;
      20'h0146b: out <= 12'h666;
      20'h0146c: out <= 12'h000;
      20'h0146d: out <= 12'h000;
      20'h0146e: out <= 12'h000;
      20'h0146f: out <= 12'h000;
      20'h01470: out <= 12'h000;
      20'h01471: out <= 12'h000;
      20'h01472: out <= 12'h000;
      20'h01473: out <= 12'h000;
      20'h01474: out <= 12'hfff;
      20'h01475: out <= 12'hbbb;
      20'h01476: out <= 12'h666;
      20'h01477: out <= 12'h666;
      20'h01478: out <= 12'h666;
      20'h01479: out <= 12'hbbb;
      20'h0147a: out <= 12'h666;
      20'h0147b: out <= 12'h666;
      20'h0147c: out <= 12'hfff;
      20'h0147d: out <= 12'hbbb;
      20'h0147e: out <= 12'h666;
      20'h0147f: out <= 12'h666;
      20'h01480: out <= 12'h666;
      20'h01481: out <= 12'hbbb;
      20'h01482: out <= 12'h666;
      20'h01483: out <= 12'h666;
      20'h01484: out <= 12'h603;
      20'h01485: out <= 12'h603;
      20'h01486: out <= 12'h603;
      20'h01487: out <= 12'h603;
      20'h01488: out <= 12'hee9;
      20'h01489: out <= 12'hf87;
      20'h0148a: out <= 12'hee9;
      20'h0148b: out <= 12'hee9;
      20'h0148c: out <= 12'hee9;
      20'h0148d: out <= 12'hb27;
      20'h0148e: out <= 12'hf87;
      20'h0148f: out <= 12'hb27;
      20'h01490: out <= 12'h000;
      20'h01491: out <= 12'h000;
      20'h01492: out <= 12'h000;
      20'h01493: out <= 12'h000;
      20'h01494: out <= 12'h000;
      20'h01495: out <= 12'h000;
      20'h01496: out <= 12'h000;
      20'h01497: out <= 12'h000;
      20'h01498: out <= 12'hee9;
      20'h01499: out <= 12'hee9;
      20'h0149a: out <= 12'hee9;
      20'h0149b: out <= 12'h000;
      20'h0149c: out <= 12'h000;
      20'h0149d: out <= 12'h000;
      20'h0149e: out <= 12'h000;
      20'h0149f: out <= 12'h000;
      20'h014a0: out <= 12'h000;
      20'h014a1: out <= 12'hee9;
      20'h014a2: out <= 12'hee9;
      20'h014a3: out <= 12'h000;
      20'h014a4: out <= 12'h000;
      20'h014a5: out <= 12'h000;
      20'h014a6: out <= 12'hee9;
      20'h014a7: out <= 12'hee9;
      20'h014a8: out <= 12'h000;
      20'h014a9: out <= 12'h000;
      20'h014aa: out <= 12'hee9;
      20'h014ab: out <= 12'hee9;
      20'h014ac: out <= 12'h000;
      20'h014ad: out <= 12'hee9;
      20'h014ae: out <= 12'hee9;
      20'h014af: out <= 12'h000;
      20'h014b0: out <= 12'h000;
      20'h014b1: out <= 12'h000;
      20'h014b2: out <= 12'h000;
      20'h014b3: out <= 12'h000;
      20'h014b4: out <= 12'hee9;
      20'h014b5: out <= 12'hee9;
      20'h014b6: out <= 12'h000;
      20'h014b7: out <= 12'h000;
      20'h014b8: out <= 12'h000;
      20'h014b9: out <= 12'h000;
      20'h014ba: out <= 12'h000;
      20'h014bb: out <= 12'h000;
      20'h014bc: out <= 12'h000;
      20'h014bd: out <= 12'h000;
      20'h014be: out <= 12'h000;
      20'h014bf: out <= 12'h000;
      20'h014c0: out <= 12'h000;
      20'h014c1: out <= 12'h000;
      20'h014c2: out <= 12'h000;
      20'h014c3: out <= 12'h000;
      20'h014c4: out <= 12'h000;
      20'h014c5: out <= 12'h000;
      20'h014c6: out <= 12'h000;
      20'h014c7: out <= 12'h000;
      20'h014c8: out <= 12'h000;
      20'h014c9: out <= 12'hfff;
      20'h014ca: out <= 12'h6af;
      20'h014cb: out <= 12'h16d;
      20'h014cc: out <= 12'h16d;
      20'h014cd: out <= 12'h16d;
      20'h014ce: out <= 12'h16d;
      20'h014cf: out <= 12'h16d;
      20'h014d0: out <= 12'h16d;
      20'h014d1: out <= 12'h16d;
      20'h014d2: out <= 12'h6af;
      20'h014d3: out <= 12'hfff;
      20'h014d4: out <= 12'h000;
      20'h014d5: out <= 12'h000;
      20'h014d6: out <= 12'h000;
      20'h014d7: out <= 12'h000;
      20'h014d8: out <= 12'h222;
      20'h014d9: out <= 12'h16d;
      20'h014da: out <= 12'h6af;
      20'h014db: out <= 12'hfff;
      20'h014dc: out <= 12'h16d;
      20'h014dd: out <= 12'h16d;
      20'h014de: out <= 12'h16d;
      20'h014df: out <= 12'h16d;
      20'h014e0: out <= 12'h16d;
      20'h014e1: out <= 12'hfff;
      20'h014e2: out <= 12'h6af;
      20'h014e3: out <= 12'h16d;
      20'h014e4: out <= 12'h222;
      20'h014e5: out <= 12'h222;
      20'h014e6: out <= 12'h222;
      20'h014e7: out <= 12'h222;
      20'h014e8: out <= 12'h000;
      20'h014e9: out <= 12'h6af;
      20'h014ea: out <= 12'h16d;
      20'h014eb: out <= 12'h6af;
      20'h014ec: out <= 12'h000;
      20'h014ed: out <= 12'h000;
      20'h014ee: out <= 12'hfff;
      20'h014ef: out <= 12'hfff;
      20'h014f0: out <= 12'hfff;
      20'h014f1: out <= 12'hfff;
      20'h014f2: out <= 12'hfff;
      20'h014f3: out <= 12'h000;
      20'h014f4: out <= 12'h000;
      20'h014f5: out <= 12'h6af;
      20'h014f6: out <= 12'h16d;
      20'h014f7: out <= 12'h6af;
      20'h014f8: out <= 12'h222;
      20'h014f9: out <= 12'h6af;
      20'h014fa: out <= 12'h16d;
      20'h014fb: out <= 12'h6af;
      20'h014fc: out <= 12'h222;
      20'h014fd: out <= 12'h222;
      20'h014fe: out <= 12'h16d;
      20'h014ff: out <= 12'h16d;
      20'h01500: out <= 12'h16d;
      20'h01501: out <= 12'h16d;
      20'h01502: out <= 12'h16d;
      20'h01503: out <= 12'h222;
      20'h01504: out <= 12'h222;
      20'h01505: out <= 12'h6af;
      20'h01506: out <= 12'h16d;
      20'h01507: out <= 12'h6af;
      20'h01508: out <= 12'h000;
      20'h01509: out <= 12'h000;
      20'h0150a: out <= 12'h000;
      20'h0150b: out <= 12'h000;
      20'h0150c: out <= 12'hfff;
      20'h0150d: out <= 12'h6af;
      20'h0150e: out <= 12'h16d;
      20'h0150f: out <= 12'h16d;
      20'h01510: out <= 12'h16d;
      20'h01511: out <= 12'h16d;
      20'h01512: out <= 12'h16d;
      20'h01513: out <= 12'h16d;
      20'h01514: out <= 12'h16d;
      20'h01515: out <= 12'h6af;
      20'h01516: out <= 12'hfff;
      20'h01517: out <= 12'h000;
      20'h01518: out <= 12'h222;
      20'h01519: out <= 12'h222;
      20'h0151a: out <= 12'h222;
      20'h0151b: out <= 12'h222;
      20'h0151c: out <= 12'h16d;
      20'h0151d: out <= 12'h6af;
      20'h0151e: out <= 12'hfff;
      20'h0151f: out <= 12'h16d;
      20'h01520: out <= 12'h16d;
      20'h01521: out <= 12'h16d;
      20'h01522: out <= 12'h16d;
      20'h01523: out <= 12'h16d;
      20'h01524: out <= 12'hfff;
      20'h01525: out <= 12'h6af;
      20'h01526: out <= 12'h16d;
      20'h01527: out <= 12'h222;
      20'h01528: out <= 12'h000;
      20'h01529: out <= 12'h6af;
      20'h0152a: out <= 12'hfff;
      20'h0152b: out <= 12'h6af;
      20'h0152c: out <= 12'h16d;
      20'h0152d: out <= 12'h16d;
      20'h0152e: out <= 12'h6af;
      20'h0152f: out <= 12'hfff;
      20'h01530: out <= 12'hfff;
      20'h01531: out <= 12'hfff;
      20'h01532: out <= 12'h6af;
      20'h01533: out <= 12'h16d;
      20'h01534: out <= 12'h16d;
      20'h01535: out <= 12'h6af;
      20'h01536: out <= 12'hfff;
      20'h01537: out <= 12'h6af;
      20'h01538: out <= 12'h222;
      20'h01539: out <= 12'h6af;
      20'h0153a: out <= 12'h16d;
      20'h0153b: out <= 12'h6af;
      20'h0153c: out <= 12'hfff;
      20'h0153d: out <= 12'hfff;
      20'h0153e: out <= 12'h6af;
      20'h0153f: out <= 12'hfff;
      20'h01540: out <= 12'hfff;
      20'h01541: out <= 12'hfff;
      20'h01542: out <= 12'h6af;
      20'h01543: out <= 12'hfff;
      20'h01544: out <= 12'hfff;
      20'h01545: out <= 12'h6af;
      20'h01546: out <= 12'h16d;
      20'h01547: out <= 12'h6af;
      20'h01548: out <= 12'h603;
      20'h01549: out <= 12'h603;
      20'h0154a: out <= 12'h603;
      20'h0154b: out <= 12'h603;
      20'h0154c: out <= 12'hfff;
      20'h0154d: out <= 12'hbbb;
      20'h0154e: out <= 12'h666;
      20'h0154f: out <= 12'hbbb;
      20'h01550: out <= 12'hfff;
      20'h01551: out <= 12'hbbb;
      20'h01552: out <= 12'h666;
      20'h01553: out <= 12'h666;
      20'h01554: out <= 12'hfff;
      20'h01555: out <= 12'hbbb;
      20'h01556: out <= 12'h666;
      20'h01557: out <= 12'hbbb;
      20'h01558: out <= 12'hfff;
      20'h01559: out <= 12'hbbb;
      20'h0155a: out <= 12'h666;
      20'h0155b: out <= 12'h666;
      20'h0155c: out <= 12'h000;
      20'h0155d: out <= 12'h000;
      20'h0155e: out <= 12'h000;
      20'h0155f: out <= 12'h000;
      20'h01560: out <= 12'h000;
      20'h01561: out <= 12'h000;
      20'h01562: out <= 12'h000;
      20'h01563: out <= 12'h000;
      20'h01564: out <= 12'hfff;
      20'h01565: out <= 12'hbbb;
      20'h01566: out <= 12'h666;
      20'h01567: out <= 12'hbbb;
      20'h01568: out <= 12'hfff;
      20'h01569: out <= 12'hbbb;
      20'h0156a: out <= 12'h666;
      20'h0156b: out <= 12'h666;
      20'h0156c: out <= 12'h000;
      20'h0156d: out <= 12'h000;
      20'h0156e: out <= 12'h000;
      20'h0156f: out <= 12'h000;
      20'h01570: out <= 12'h000;
      20'h01571: out <= 12'h000;
      20'h01572: out <= 12'h000;
      20'h01573: out <= 12'h000;
      20'h01574: out <= 12'h000;
      20'h01575: out <= 12'h000;
      20'h01576: out <= 12'h000;
      20'h01577: out <= 12'h000;
      20'h01578: out <= 12'h000;
      20'h01579: out <= 12'h000;
      20'h0157a: out <= 12'h000;
      20'h0157b: out <= 12'h000;
      20'h0157c: out <= 12'hfff;
      20'h0157d: out <= 12'hbbb;
      20'h0157e: out <= 12'h666;
      20'h0157f: out <= 12'hbbb;
      20'h01580: out <= 12'hfff;
      20'h01581: out <= 12'hbbb;
      20'h01582: out <= 12'h666;
      20'h01583: out <= 12'h666;
      20'h01584: out <= 12'h000;
      20'h01585: out <= 12'h000;
      20'h01586: out <= 12'h000;
      20'h01587: out <= 12'h000;
      20'h01588: out <= 12'h000;
      20'h01589: out <= 12'h000;
      20'h0158a: out <= 12'h000;
      20'h0158b: out <= 12'h000;
      20'h0158c: out <= 12'hfff;
      20'h0158d: out <= 12'hbbb;
      20'h0158e: out <= 12'h666;
      20'h0158f: out <= 12'hbbb;
      20'h01590: out <= 12'hfff;
      20'h01591: out <= 12'hbbb;
      20'h01592: out <= 12'h666;
      20'h01593: out <= 12'h666;
      20'h01594: out <= 12'hfff;
      20'h01595: out <= 12'hbbb;
      20'h01596: out <= 12'h666;
      20'h01597: out <= 12'hbbb;
      20'h01598: out <= 12'hfff;
      20'h01599: out <= 12'hbbb;
      20'h0159a: out <= 12'h666;
      20'h0159b: out <= 12'h666;
      20'h0159c: out <= 12'h603;
      20'h0159d: out <= 12'h603;
      20'h0159e: out <= 12'h603;
      20'h0159f: out <= 12'h603;
      20'h015a0: out <= 12'hee9;
      20'h015a1: out <= 12'hf87;
      20'h015a2: out <= 12'hee9;
      20'h015a3: out <= 12'hf87;
      20'h015a4: out <= 12'hf87;
      20'h015a5: out <= 12'hb27;
      20'h015a6: out <= 12'hf87;
      20'h015a7: out <= 12'hb27;
      20'h015a8: out <= 12'h000;
      20'h015a9: out <= 12'h000;
      20'h015aa: out <= 12'h000;
      20'h015ab: out <= 12'h000;
      20'h015ac: out <= 12'h000;
      20'h015ad: out <= 12'h000;
      20'h015ae: out <= 12'h000;
      20'h015af: out <= 12'h000;
      20'h015b0: out <= 12'h000;
      20'h015b1: out <= 12'hee9;
      20'h015b2: out <= 12'hee9;
      20'h015b3: out <= 12'hee9;
      20'h015b4: out <= 12'hee9;
      20'h015b5: out <= 12'h000;
      20'h015b6: out <= 12'h000;
      20'h015b7: out <= 12'h000;
      20'h015b8: out <= 12'h000;
      20'h015b9: out <= 12'hee9;
      20'h015ba: out <= 12'hee9;
      20'h015bb: out <= 12'h000;
      20'h015bc: out <= 12'h000;
      20'h015bd: out <= 12'h000;
      20'h015be: out <= 12'hee9;
      20'h015bf: out <= 12'hee9;
      20'h015c0: out <= 12'h000;
      20'h015c1: out <= 12'h000;
      20'h015c2: out <= 12'hee9;
      20'h015c3: out <= 12'hee9;
      20'h015c4: out <= 12'h000;
      20'h015c5: out <= 12'hee9;
      20'h015c6: out <= 12'hee9;
      20'h015c7: out <= 12'h000;
      20'h015c8: out <= 12'h000;
      20'h015c9: out <= 12'h000;
      20'h015ca: out <= 12'h000;
      20'h015cb: out <= 12'h000;
      20'h015cc: out <= 12'hee9;
      20'h015cd: out <= 12'hee9;
      20'h015ce: out <= 12'hee9;
      20'h015cf: out <= 12'hee9;
      20'h015d0: out <= 12'h000;
      20'h015d1: out <= 12'h000;
      20'h015d2: out <= 12'h000;
      20'h015d3: out <= 12'h000;
      20'h015d4: out <= 12'h000;
      20'h015d5: out <= 12'h000;
      20'h015d6: out <= 12'h000;
      20'h015d7: out <= 12'h000;
      20'h015d8: out <= 12'h000;
      20'h015d9: out <= 12'h000;
      20'h015da: out <= 12'h000;
      20'h015db: out <= 12'h000;
      20'h015dc: out <= 12'h000;
      20'h015dd: out <= 12'h000;
      20'h015de: out <= 12'h000;
      20'h015df: out <= 12'h000;
      20'h015e0: out <= 12'h000;
      20'h015e1: out <= 12'hfff;
      20'h015e2: out <= 12'h6af;
      20'h015e3: out <= 12'h16d;
      20'h015e4: out <= 12'h6af;
      20'h015e5: out <= 12'h16d;
      20'h015e6: out <= 12'h16d;
      20'h015e7: out <= 12'h16d;
      20'h015e8: out <= 12'h16d;
      20'h015e9: out <= 12'h16d;
      20'h015ea: out <= 12'h6af;
      20'h015eb: out <= 12'hfff;
      20'h015ec: out <= 12'h000;
      20'h015ed: out <= 12'h000;
      20'h015ee: out <= 12'h000;
      20'h015ef: out <= 12'h000;
      20'h015f0: out <= 12'h222;
      20'h015f1: out <= 12'h16d;
      20'h015f2: out <= 12'h6af;
      20'h015f3: out <= 12'hfff;
      20'h015f4: out <= 12'h6af;
      20'h015f5: out <= 12'h16d;
      20'h015f6: out <= 12'h16d;
      20'h015f7: out <= 12'h16d;
      20'h015f8: out <= 12'h16d;
      20'h015f9: out <= 12'hfff;
      20'h015fa: out <= 12'h6af;
      20'h015fb: out <= 12'h16d;
      20'h015fc: out <= 12'h222;
      20'h015fd: out <= 12'h222;
      20'h015fe: out <= 12'h222;
      20'h015ff: out <= 12'h222;
      20'h01600: out <= 12'h000;
      20'h01601: out <= 12'hfff;
      20'h01602: out <= 12'hfff;
      20'h01603: out <= 12'hfff;
      20'h01604: out <= 12'hfff;
      20'h01605: out <= 12'hfff;
      20'h01606: out <= 12'h6af;
      20'h01607: out <= 12'h6af;
      20'h01608: out <= 12'h6af;
      20'h01609: out <= 12'h6af;
      20'h0160a: out <= 12'h6af;
      20'h0160b: out <= 12'hfff;
      20'h0160c: out <= 12'hfff;
      20'h0160d: out <= 12'hfff;
      20'h0160e: out <= 12'hfff;
      20'h0160f: out <= 12'hfff;
      20'h01610: out <= 12'h222;
      20'h01611: out <= 12'hfff;
      20'h01612: out <= 12'hfff;
      20'h01613: out <= 12'hfff;
      20'h01614: out <= 12'h16d;
      20'h01615: out <= 12'h16d;
      20'h01616: out <= 12'h6af;
      20'h01617: out <= 12'h6af;
      20'h01618: out <= 12'h6af;
      20'h01619: out <= 12'h6af;
      20'h0161a: out <= 12'h6af;
      20'h0161b: out <= 12'h16d;
      20'h0161c: out <= 12'h16d;
      20'h0161d: out <= 12'hfff;
      20'h0161e: out <= 12'hfff;
      20'h0161f: out <= 12'hfff;
      20'h01620: out <= 12'h000;
      20'h01621: out <= 12'h000;
      20'h01622: out <= 12'h000;
      20'h01623: out <= 12'h000;
      20'h01624: out <= 12'hfff;
      20'h01625: out <= 12'h6af;
      20'h01626: out <= 12'h16d;
      20'h01627: out <= 12'h16d;
      20'h01628: out <= 12'h16d;
      20'h01629: out <= 12'h16d;
      20'h0162a: out <= 12'h16d;
      20'h0162b: out <= 12'h6af;
      20'h0162c: out <= 12'h16d;
      20'h0162d: out <= 12'h6af;
      20'h0162e: out <= 12'hfff;
      20'h0162f: out <= 12'h000;
      20'h01630: out <= 12'h222;
      20'h01631: out <= 12'h222;
      20'h01632: out <= 12'h222;
      20'h01633: out <= 12'h222;
      20'h01634: out <= 12'h16d;
      20'h01635: out <= 12'h6af;
      20'h01636: out <= 12'hfff;
      20'h01637: out <= 12'h16d;
      20'h01638: out <= 12'h16d;
      20'h01639: out <= 12'h16d;
      20'h0163a: out <= 12'h16d;
      20'h0163b: out <= 12'h6af;
      20'h0163c: out <= 12'hfff;
      20'h0163d: out <= 12'h6af;
      20'h0163e: out <= 12'h16d;
      20'h0163f: out <= 12'h222;
      20'h01640: out <= 12'h000;
      20'h01641: out <= 12'hfff;
      20'h01642: out <= 12'h6af;
      20'h01643: out <= 12'h16d;
      20'h01644: out <= 12'h16d;
      20'h01645: out <= 12'h6af;
      20'h01646: out <= 12'h16d;
      20'h01647: out <= 12'h16d;
      20'h01648: out <= 12'h16d;
      20'h01649: out <= 12'h16d;
      20'h0164a: out <= 12'h16d;
      20'h0164b: out <= 12'h6af;
      20'h0164c: out <= 12'h16d;
      20'h0164d: out <= 12'h16d;
      20'h0164e: out <= 12'h6af;
      20'h0164f: out <= 12'hfff;
      20'h01650: out <= 12'h222;
      20'h01651: out <= 12'h16d;
      20'h01652: out <= 12'h6af;
      20'h01653: out <= 12'hfff;
      20'h01654: out <= 12'h16d;
      20'h01655: out <= 12'h6af;
      20'h01656: out <= 12'h16d;
      20'h01657: out <= 12'h16d;
      20'h01658: out <= 12'h16d;
      20'h01659: out <= 12'h16d;
      20'h0165a: out <= 12'h16d;
      20'h0165b: out <= 12'h6af;
      20'h0165c: out <= 12'h16d;
      20'h0165d: out <= 12'hfff;
      20'h0165e: out <= 12'h6af;
      20'h0165f: out <= 12'h16d;
      20'h01660: out <= 12'h603;
      20'h01661: out <= 12'h603;
      20'h01662: out <= 12'h603;
      20'h01663: out <= 12'h603;
      20'h01664: out <= 12'hfff;
      20'h01665: out <= 12'hbbb;
      20'h01666: out <= 12'h666;
      20'h01667: out <= 12'hfff;
      20'h01668: out <= 12'hfff;
      20'h01669: out <= 12'hbbb;
      20'h0166a: out <= 12'h666;
      20'h0166b: out <= 12'h666;
      20'h0166c: out <= 12'hfff;
      20'h0166d: out <= 12'hbbb;
      20'h0166e: out <= 12'h666;
      20'h0166f: out <= 12'hfff;
      20'h01670: out <= 12'hfff;
      20'h01671: out <= 12'hbbb;
      20'h01672: out <= 12'h666;
      20'h01673: out <= 12'h666;
      20'h01674: out <= 12'h000;
      20'h01675: out <= 12'h000;
      20'h01676: out <= 12'h000;
      20'h01677: out <= 12'h000;
      20'h01678: out <= 12'h000;
      20'h01679: out <= 12'h000;
      20'h0167a: out <= 12'h000;
      20'h0167b: out <= 12'h000;
      20'h0167c: out <= 12'hfff;
      20'h0167d: out <= 12'hbbb;
      20'h0167e: out <= 12'h666;
      20'h0167f: out <= 12'hfff;
      20'h01680: out <= 12'hfff;
      20'h01681: out <= 12'hbbb;
      20'h01682: out <= 12'h666;
      20'h01683: out <= 12'h666;
      20'h01684: out <= 12'h000;
      20'h01685: out <= 12'h000;
      20'h01686: out <= 12'h000;
      20'h01687: out <= 12'h000;
      20'h01688: out <= 12'h000;
      20'h01689: out <= 12'h000;
      20'h0168a: out <= 12'h000;
      20'h0168b: out <= 12'h000;
      20'h0168c: out <= 12'h000;
      20'h0168d: out <= 12'h000;
      20'h0168e: out <= 12'h000;
      20'h0168f: out <= 12'h000;
      20'h01690: out <= 12'h000;
      20'h01691: out <= 12'h000;
      20'h01692: out <= 12'h000;
      20'h01693: out <= 12'h000;
      20'h01694: out <= 12'hfff;
      20'h01695: out <= 12'hbbb;
      20'h01696: out <= 12'h666;
      20'h01697: out <= 12'hfff;
      20'h01698: out <= 12'hfff;
      20'h01699: out <= 12'hbbb;
      20'h0169a: out <= 12'h666;
      20'h0169b: out <= 12'h666;
      20'h0169c: out <= 12'h000;
      20'h0169d: out <= 12'h000;
      20'h0169e: out <= 12'h000;
      20'h0169f: out <= 12'h000;
      20'h016a0: out <= 12'h000;
      20'h016a1: out <= 12'h000;
      20'h016a2: out <= 12'h000;
      20'h016a3: out <= 12'h000;
      20'h016a4: out <= 12'hfff;
      20'h016a5: out <= 12'hbbb;
      20'h016a6: out <= 12'h666;
      20'h016a7: out <= 12'hfff;
      20'h016a8: out <= 12'hfff;
      20'h016a9: out <= 12'hbbb;
      20'h016aa: out <= 12'h666;
      20'h016ab: out <= 12'h666;
      20'h016ac: out <= 12'hfff;
      20'h016ad: out <= 12'hbbb;
      20'h016ae: out <= 12'h666;
      20'h016af: out <= 12'hfff;
      20'h016b0: out <= 12'hfff;
      20'h016b1: out <= 12'hbbb;
      20'h016b2: out <= 12'h666;
      20'h016b3: out <= 12'h666;
      20'h016b4: out <= 12'h603;
      20'h016b5: out <= 12'h603;
      20'h016b6: out <= 12'h603;
      20'h016b7: out <= 12'h603;
      20'h016b8: out <= 12'hee9;
      20'h016b9: out <= 12'hf87;
      20'h016ba: out <= 12'hee9;
      20'h016bb: out <= 12'hf87;
      20'h016bc: out <= 12'hf87;
      20'h016bd: out <= 12'hb27;
      20'h016be: out <= 12'hf87;
      20'h016bf: out <= 12'hb27;
      20'h016c0: out <= 12'h000;
      20'h016c1: out <= 12'h000;
      20'h016c2: out <= 12'h000;
      20'h016c3: out <= 12'h000;
      20'h016c4: out <= 12'h000;
      20'h016c5: out <= 12'h000;
      20'h016c6: out <= 12'h000;
      20'h016c7: out <= 12'h000;
      20'h016c8: out <= 12'h000;
      20'h016c9: out <= 12'h000;
      20'h016ca: out <= 12'h000;
      20'h016cb: out <= 12'hee9;
      20'h016cc: out <= 12'hee9;
      20'h016cd: out <= 12'hee9;
      20'h016ce: out <= 12'h000;
      20'h016cf: out <= 12'h000;
      20'h016d0: out <= 12'h000;
      20'h016d1: out <= 12'hee9;
      20'h016d2: out <= 12'hee9;
      20'h016d3: out <= 12'h000;
      20'h016d4: out <= 12'h000;
      20'h016d5: out <= 12'h000;
      20'h016d6: out <= 12'hee9;
      20'h016d7: out <= 12'hee9;
      20'h016d8: out <= 12'hee9;
      20'h016d9: out <= 12'hee9;
      20'h016da: out <= 12'hee9;
      20'h016db: out <= 12'hee9;
      20'h016dc: out <= 12'h000;
      20'h016dd: out <= 12'hee9;
      20'h016de: out <= 12'hee9;
      20'h016df: out <= 12'h000;
      20'h016e0: out <= 12'hee9;
      20'h016e1: out <= 12'hee9;
      20'h016e2: out <= 12'hee9;
      20'h016e3: out <= 12'h000;
      20'h016e4: out <= 12'hee9;
      20'h016e5: out <= 12'hee9;
      20'h016e6: out <= 12'h000;
      20'h016e7: out <= 12'h000;
      20'h016e8: out <= 12'h000;
      20'h016e9: out <= 12'h000;
      20'h016ea: out <= 12'h000;
      20'h016eb: out <= 12'h000;
      20'h016ec: out <= 12'h000;
      20'h016ed: out <= 12'h000;
      20'h016ee: out <= 12'h000;
      20'h016ef: out <= 12'h000;
      20'h016f0: out <= 12'h000;
      20'h016f1: out <= 12'h000;
      20'h016f2: out <= 12'h000;
      20'h016f3: out <= 12'h000;
      20'h016f4: out <= 12'h000;
      20'h016f5: out <= 12'h000;
      20'h016f6: out <= 12'h000;
      20'h016f7: out <= 12'h000;
      20'h016f8: out <= 12'hfff;
      20'h016f9: out <= 12'h6af;
      20'h016fa: out <= 12'h16d;
      20'h016fb: out <= 12'h6af;
      20'h016fc: out <= 12'h16d;
      20'h016fd: out <= 12'h16d;
      20'h016fe: out <= 12'h6af;
      20'h016ff: out <= 12'h6af;
      20'h01700: out <= 12'h16d;
      20'h01701: out <= 12'h16d;
      20'h01702: out <= 12'h16d;
      20'h01703: out <= 12'h6af;
      20'h01704: out <= 12'hfff;
      20'h01705: out <= 12'h000;
      20'h01706: out <= 12'h000;
      20'h01707: out <= 12'h000;
      20'h01708: out <= 12'h16d;
      20'h01709: out <= 12'h6af;
      20'h0170a: out <= 12'hfff;
      20'h0170b: out <= 12'h6af;
      20'h0170c: out <= 12'h16d;
      20'h0170d: out <= 12'h16d;
      20'h0170e: out <= 12'h6af;
      20'h0170f: out <= 12'h6af;
      20'h01710: out <= 12'h16d;
      20'h01711: out <= 12'h16d;
      20'h01712: out <= 12'hfff;
      20'h01713: out <= 12'h6af;
      20'h01714: out <= 12'h16d;
      20'h01715: out <= 12'h222;
      20'h01716: out <= 12'h222;
      20'h01717: out <= 12'h222;
      20'h01718: out <= 12'h000;
      20'h01719: out <= 12'h6af;
      20'h0171a: out <= 12'h16d;
      20'h0171b: out <= 12'hfff;
      20'h0171c: out <= 12'h6af;
      20'h0171d: out <= 12'h6af;
      20'h0171e: out <= 12'h16d;
      20'h0171f: out <= 12'h16d;
      20'h01720: out <= 12'h16d;
      20'h01721: out <= 12'h16d;
      20'h01722: out <= 12'h16d;
      20'h01723: out <= 12'h6af;
      20'h01724: out <= 12'h6af;
      20'h01725: out <= 12'hfff;
      20'h01726: out <= 12'h16d;
      20'h01727: out <= 12'h6af;
      20'h01728: out <= 12'h222;
      20'h01729: out <= 12'h6af;
      20'h0172a: out <= 12'h16d;
      20'h0172b: out <= 12'h16d;
      20'h0172c: out <= 12'h6af;
      20'h0172d: out <= 12'h6af;
      20'h0172e: out <= 12'hfff;
      20'h0172f: out <= 12'hfff;
      20'h01730: out <= 12'hfff;
      20'h01731: out <= 12'hfff;
      20'h01732: out <= 12'hfff;
      20'h01733: out <= 12'h6af;
      20'h01734: out <= 12'h6af;
      20'h01735: out <= 12'h16d;
      20'h01736: out <= 12'h16d;
      20'h01737: out <= 12'h6af;
      20'h01738: out <= 12'h000;
      20'h01739: out <= 12'h000;
      20'h0173a: out <= 12'h000;
      20'h0173b: out <= 12'hfff;
      20'h0173c: out <= 12'h6af;
      20'h0173d: out <= 12'h16d;
      20'h0173e: out <= 12'h16d;
      20'h0173f: out <= 12'h16d;
      20'h01740: out <= 12'h6af;
      20'h01741: out <= 12'h6af;
      20'h01742: out <= 12'h16d;
      20'h01743: out <= 12'h16d;
      20'h01744: out <= 12'h6af;
      20'h01745: out <= 12'h16d;
      20'h01746: out <= 12'h6af;
      20'h01747: out <= 12'hfff;
      20'h01748: out <= 12'h222;
      20'h01749: out <= 12'h222;
      20'h0174a: out <= 12'h222;
      20'h0174b: out <= 12'h16d;
      20'h0174c: out <= 12'h6af;
      20'h0174d: out <= 12'hfff;
      20'h0174e: out <= 12'h16d;
      20'h0174f: out <= 12'h16d;
      20'h01750: out <= 12'h6af;
      20'h01751: out <= 12'h6af;
      20'h01752: out <= 12'h16d;
      20'h01753: out <= 12'h16d;
      20'h01754: out <= 12'h6af;
      20'h01755: out <= 12'hfff;
      20'h01756: out <= 12'h6af;
      20'h01757: out <= 12'h16d;
      20'h01758: out <= 12'h000;
      20'h01759: out <= 12'hfff;
      20'h0175a: out <= 12'h6af;
      20'h0175b: out <= 12'h16d;
      20'h0175c: out <= 12'h16d;
      20'h0175d: out <= 12'h16d;
      20'h0175e: out <= 12'h16d;
      20'h0175f: out <= 12'h6af;
      20'h01760: out <= 12'hfff;
      20'h01761: out <= 12'h6af;
      20'h01762: out <= 12'h16d;
      20'h01763: out <= 12'h16d;
      20'h01764: out <= 12'h16d;
      20'h01765: out <= 12'h16d;
      20'h01766: out <= 12'h6af;
      20'h01767: out <= 12'hfff;
      20'h01768: out <= 12'h222;
      20'h01769: out <= 12'h16d;
      20'h0176a: out <= 12'h6af;
      20'h0176b: out <= 12'hfff;
      20'h0176c: out <= 12'h16d;
      20'h0176d: out <= 12'h16d;
      20'h0176e: out <= 12'h16d;
      20'h0176f: out <= 12'h6af;
      20'h01770: out <= 12'hfff;
      20'h01771: out <= 12'h6af;
      20'h01772: out <= 12'h16d;
      20'h01773: out <= 12'h16d;
      20'h01774: out <= 12'h16d;
      20'h01775: out <= 12'hfff;
      20'h01776: out <= 12'h6af;
      20'h01777: out <= 12'h16d;
      20'h01778: out <= 12'h603;
      20'h01779: out <= 12'h603;
      20'h0177a: out <= 12'h603;
      20'h0177b: out <= 12'h603;
      20'h0177c: out <= 12'hfff;
      20'h0177d: out <= 12'hbbb;
      20'h0177e: out <= 12'hbbb;
      20'h0177f: out <= 12'hbbb;
      20'h01780: out <= 12'hbbb;
      20'h01781: out <= 12'hbbb;
      20'h01782: out <= 12'h666;
      20'h01783: out <= 12'h666;
      20'h01784: out <= 12'hfff;
      20'h01785: out <= 12'hbbb;
      20'h01786: out <= 12'hbbb;
      20'h01787: out <= 12'hbbb;
      20'h01788: out <= 12'hbbb;
      20'h01789: out <= 12'hbbb;
      20'h0178a: out <= 12'h666;
      20'h0178b: out <= 12'h666;
      20'h0178c: out <= 12'h000;
      20'h0178d: out <= 12'h000;
      20'h0178e: out <= 12'h000;
      20'h0178f: out <= 12'h000;
      20'h01790: out <= 12'h000;
      20'h01791: out <= 12'h000;
      20'h01792: out <= 12'h000;
      20'h01793: out <= 12'h000;
      20'h01794: out <= 12'hfff;
      20'h01795: out <= 12'hbbb;
      20'h01796: out <= 12'hbbb;
      20'h01797: out <= 12'hbbb;
      20'h01798: out <= 12'hbbb;
      20'h01799: out <= 12'hbbb;
      20'h0179a: out <= 12'h666;
      20'h0179b: out <= 12'h666;
      20'h0179c: out <= 12'h000;
      20'h0179d: out <= 12'h000;
      20'h0179e: out <= 12'h000;
      20'h0179f: out <= 12'h000;
      20'h017a0: out <= 12'h000;
      20'h017a1: out <= 12'h000;
      20'h017a2: out <= 12'h000;
      20'h017a3: out <= 12'h000;
      20'h017a4: out <= 12'h000;
      20'h017a5: out <= 12'h000;
      20'h017a6: out <= 12'h000;
      20'h017a7: out <= 12'h000;
      20'h017a8: out <= 12'h000;
      20'h017a9: out <= 12'h000;
      20'h017aa: out <= 12'h000;
      20'h017ab: out <= 12'h000;
      20'h017ac: out <= 12'hfff;
      20'h017ad: out <= 12'hbbb;
      20'h017ae: out <= 12'hbbb;
      20'h017af: out <= 12'hbbb;
      20'h017b0: out <= 12'hbbb;
      20'h017b1: out <= 12'hbbb;
      20'h017b2: out <= 12'h666;
      20'h017b3: out <= 12'h666;
      20'h017b4: out <= 12'h000;
      20'h017b5: out <= 12'h000;
      20'h017b6: out <= 12'h000;
      20'h017b7: out <= 12'h000;
      20'h017b8: out <= 12'h000;
      20'h017b9: out <= 12'h000;
      20'h017ba: out <= 12'h000;
      20'h017bb: out <= 12'h000;
      20'h017bc: out <= 12'hfff;
      20'h017bd: out <= 12'hbbb;
      20'h017be: out <= 12'hbbb;
      20'h017bf: out <= 12'hbbb;
      20'h017c0: out <= 12'hbbb;
      20'h017c1: out <= 12'hbbb;
      20'h017c2: out <= 12'h666;
      20'h017c3: out <= 12'h666;
      20'h017c4: out <= 12'hfff;
      20'h017c5: out <= 12'hbbb;
      20'h017c6: out <= 12'hbbb;
      20'h017c7: out <= 12'hbbb;
      20'h017c8: out <= 12'hbbb;
      20'h017c9: out <= 12'hbbb;
      20'h017ca: out <= 12'h666;
      20'h017cb: out <= 12'h666;
      20'h017cc: out <= 12'h603;
      20'h017cd: out <= 12'h603;
      20'h017ce: out <= 12'h603;
      20'h017cf: out <= 12'h603;
      20'h017d0: out <= 12'hee9;
      20'h017d1: out <= 12'hf87;
      20'h017d2: out <= 12'hee9;
      20'h017d3: out <= 12'hb27;
      20'h017d4: out <= 12'hb27;
      20'h017d5: out <= 12'hb27;
      20'h017d6: out <= 12'hf87;
      20'h017d7: out <= 12'hb27;
      20'h017d8: out <= 12'h000;
      20'h017d9: out <= 12'h000;
      20'h017da: out <= 12'h000;
      20'h017db: out <= 12'h000;
      20'h017dc: out <= 12'h000;
      20'h017dd: out <= 12'h000;
      20'h017de: out <= 12'h000;
      20'h017df: out <= 12'h000;
      20'h017e0: out <= 12'hee9;
      20'h017e1: out <= 12'hee9;
      20'h017e2: out <= 12'h000;
      20'h017e3: out <= 12'h000;
      20'h017e4: out <= 12'hee9;
      20'h017e5: out <= 12'hee9;
      20'h017e6: out <= 12'h000;
      20'h017e7: out <= 12'h000;
      20'h017e8: out <= 12'h000;
      20'h017e9: out <= 12'hee9;
      20'h017ea: out <= 12'hee9;
      20'h017eb: out <= 12'h000;
      20'h017ec: out <= 12'h000;
      20'h017ed: out <= 12'h000;
      20'h017ee: out <= 12'hee9;
      20'h017ef: out <= 12'hee9;
      20'h017f0: out <= 12'h000;
      20'h017f1: out <= 12'h000;
      20'h017f2: out <= 12'hee9;
      20'h017f3: out <= 12'hee9;
      20'h017f4: out <= 12'h000;
      20'h017f5: out <= 12'hee9;
      20'h017f6: out <= 12'hee9;
      20'h017f7: out <= 12'h000;
      20'h017f8: out <= 12'h000;
      20'h017f9: out <= 12'hee9;
      20'h017fa: out <= 12'hee9;
      20'h017fb: out <= 12'h000;
      20'h017fc: out <= 12'hee9;
      20'h017fd: out <= 12'hee9;
      20'h017fe: out <= 12'h000;
      20'h017ff: out <= 12'h000;
      20'h01800: out <= 12'h000;
      20'h01801: out <= 12'h000;
      20'h01802: out <= 12'h000;
      20'h01803: out <= 12'h000;
      20'h01804: out <= 12'h000;
      20'h01805: out <= 12'h000;
      20'h01806: out <= 12'h000;
      20'h01807: out <= 12'h000;
      20'h01808: out <= 12'h000;
      20'h01809: out <= 12'h000;
      20'h0180a: out <= 12'h000;
      20'h0180b: out <= 12'h000;
      20'h0180c: out <= 12'h000;
      20'h0180d: out <= 12'h000;
      20'h0180e: out <= 12'h000;
      20'h0180f: out <= 12'h000;
      20'h01810: out <= 12'hfff;
      20'h01811: out <= 12'h6af;
      20'h01812: out <= 12'h16d;
      20'h01813: out <= 12'hfff;
      20'h01814: out <= 12'h16d;
      20'h01815: out <= 12'h6af;
      20'h01816: out <= 12'hfff;
      20'h01817: out <= 12'hfff;
      20'h01818: out <= 12'h6af;
      20'h01819: out <= 12'h16d;
      20'h0181a: out <= 12'h16d;
      20'h0181b: out <= 12'h6af;
      20'h0181c: out <= 12'hfff;
      20'h0181d: out <= 12'h16d;
      20'h0181e: out <= 12'h16d;
      20'h0181f: out <= 12'h6af;
      20'h01820: out <= 12'h16d;
      20'h01821: out <= 12'h6af;
      20'h01822: out <= 12'hfff;
      20'h01823: out <= 12'hfff;
      20'h01824: out <= 12'h16d;
      20'h01825: out <= 12'h6af;
      20'h01826: out <= 12'hfff;
      20'h01827: out <= 12'hfff;
      20'h01828: out <= 12'h6af;
      20'h01829: out <= 12'h16d;
      20'h0182a: out <= 12'hfff;
      20'h0182b: out <= 12'h6af;
      20'h0182c: out <= 12'h16d;
      20'h0182d: out <= 12'h16d;
      20'h0182e: out <= 12'h16d;
      20'h0182f: out <= 12'h6af;
      20'h01830: out <= 12'h000;
      20'h01831: out <= 12'h6af;
      20'h01832: out <= 12'hfff;
      20'h01833: out <= 12'h6af;
      20'h01834: out <= 12'h16d;
      20'h01835: out <= 12'h16d;
      20'h01836: out <= 12'h16d;
      20'h01837: out <= 12'h16d;
      20'h01838: out <= 12'h16d;
      20'h01839: out <= 12'h16d;
      20'h0183a: out <= 12'h16d;
      20'h0183b: out <= 12'h16d;
      20'h0183c: out <= 12'h16d;
      20'h0183d: out <= 12'h6af;
      20'h0183e: out <= 12'hfff;
      20'h0183f: out <= 12'h6af;
      20'h01840: out <= 12'h222;
      20'h01841: out <= 12'h6af;
      20'h01842: out <= 12'h16d;
      20'h01843: out <= 12'h6af;
      20'h01844: out <= 12'hfff;
      20'h01845: out <= 12'hfff;
      20'h01846: out <= 12'h16d;
      20'h01847: out <= 12'h16d;
      20'h01848: out <= 12'h16d;
      20'h01849: out <= 12'h16d;
      20'h0184a: out <= 12'h16d;
      20'h0184b: out <= 12'hfff;
      20'h0184c: out <= 12'hfff;
      20'h0184d: out <= 12'h6af;
      20'h0184e: out <= 12'h16d;
      20'h0184f: out <= 12'h6af;
      20'h01850: out <= 12'h6af;
      20'h01851: out <= 12'h16d;
      20'h01852: out <= 12'h16d;
      20'h01853: out <= 12'hfff;
      20'h01854: out <= 12'h6af;
      20'h01855: out <= 12'h16d;
      20'h01856: out <= 12'h16d;
      20'h01857: out <= 12'h6af;
      20'h01858: out <= 12'hfff;
      20'h01859: out <= 12'hfff;
      20'h0185a: out <= 12'h6af;
      20'h0185b: out <= 12'h16d;
      20'h0185c: out <= 12'hfff;
      20'h0185d: out <= 12'h16d;
      20'h0185e: out <= 12'h6af;
      20'h0185f: out <= 12'hfff;
      20'h01860: out <= 12'h6af;
      20'h01861: out <= 12'h16d;
      20'h01862: out <= 12'h16d;
      20'h01863: out <= 12'h16d;
      20'h01864: out <= 12'h6af;
      20'h01865: out <= 12'hfff;
      20'h01866: out <= 12'h16d;
      20'h01867: out <= 12'h6af;
      20'h01868: out <= 12'hfff;
      20'h01869: out <= 12'hfff;
      20'h0186a: out <= 12'h6af;
      20'h0186b: out <= 12'h16d;
      20'h0186c: out <= 12'hfff;
      20'h0186d: out <= 12'hfff;
      20'h0186e: out <= 12'h6af;
      20'h0186f: out <= 12'h16d;
      20'h01870: out <= 12'h000;
      20'h01871: out <= 12'hfff;
      20'h01872: out <= 12'h6af;
      20'h01873: out <= 12'h16d;
      20'h01874: out <= 12'h16d;
      20'h01875: out <= 12'h16d;
      20'h01876: out <= 12'h6af;
      20'h01877: out <= 12'hfff;
      20'h01878: out <= 12'hfff;
      20'h01879: out <= 12'hfff;
      20'h0187a: out <= 12'h6af;
      20'h0187b: out <= 12'h16d;
      20'h0187c: out <= 12'h16d;
      20'h0187d: out <= 12'h16d;
      20'h0187e: out <= 12'h6af;
      20'h0187f: out <= 12'hfff;
      20'h01880: out <= 12'h222;
      20'h01881: out <= 12'h16d;
      20'h01882: out <= 12'h6af;
      20'h01883: out <= 12'hfff;
      20'h01884: out <= 12'h16d;
      20'h01885: out <= 12'h16d;
      20'h01886: out <= 12'h6af;
      20'h01887: out <= 12'hfff;
      20'h01888: out <= 12'hfff;
      20'h01889: out <= 12'hfff;
      20'h0188a: out <= 12'h6af;
      20'h0188b: out <= 12'h16d;
      20'h0188c: out <= 12'h16d;
      20'h0188d: out <= 12'hfff;
      20'h0188e: out <= 12'h6af;
      20'h0188f: out <= 12'h16d;
      20'h01890: out <= 12'h603;
      20'h01891: out <= 12'h603;
      20'h01892: out <= 12'h603;
      20'h01893: out <= 12'h603;
      20'h01894: out <= 12'hfff;
      20'h01895: out <= 12'h666;
      20'h01896: out <= 12'h666;
      20'h01897: out <= 12'h666;
      20'h01898: out <= 12'h666;
      20'h01899: out <= 12'h666;
      20'h0189a: out <= 12'h666;
      20'h0189b: out <= 12'h666;
      20'h0189c: out <= 12'hfff;
      20'h0189d: out <= 12'h666;
      20'h0189e: out <= 12'h666;
      20'h0189f: out <= 12'h666;
      20'h018a0: out <= 12'h666;
      20'h018a1: out <= 12'h666;
      20'h018a2: out <= 12'h666;
      20'h018a3: out <= 12'h666;
      20'h018a4: out <= 12'h000;
      20'h018a5: out <= 12'h000;
      20'h018a6: out <= 12'h000;
      20'h018a7: out <= 12'h000;
      20'h018a8: out <= 12'h000;
      20'h018a9: out <= 12'h000;
      20'h018aa: out <= 12'h000;
      20'h018ab: out <= 12'h000;
      20'h018ac: out <= 12'hfff;
      20'h018ad: out <= 12'h666;
      20'h018ae: out <= 12'h666;
      20'h018af: out <= 12'h666;
      20'h018b0: out <= 12'h666;
      20'h018b1: out <= 12'h666;
      20'h018b2: out <= 12'h666;
      20'h018b3: out <= 12'h666;
      20'h018b4: out <= 12'h000;
      20'h018b5: out <= 12'h000;
      20'h018b6: out <= 12'h000;
      20'h018b7: out <= 12'h000;
      20'h018b8: out <= 12'h000;
      20'h018b9: out <= 12'h000;
      20'h018ba: out <= 12'h000;
      20'h018bb: out <= 12'h000;
      20'h018bc: out <= 12'h000;
      20'h018bd: out <= 12'h000;
      20'h018be: out <= 12'h000;
      20'h018bf: out <= 12'h000;
      20'h018c0: out <= 12'h000;
      20'h018c1: out <= 12'h000;
      20'h018c2: out <= 12'h000;
      20'h018c3: out <= 12'h000;
      20'h018c4: out <= 12'hfff;
      20'h018c5: out <= 12'h666;
      20'h018c6: out <= 12'h666;
      20'h018c7: out <= 12'h666;
      20'h018c8: out <= 12'h666;
      20'h018c9: out <= 12'h666;
      20'h018ca: out <= 12'h666;
      20'h018cb: out <= 12'h666;
      20'h018cc: out <= 12'h000;
      20'h018cd: out <= 12'h000;
      20'h018ce: out <= 12'h000;
      20'h018cf: out <= 12'h000;
      20'h018d0: out <= 12'h000;
      20'h018d1: out <= 12'h000;
      20'h018d2: out <= 12'h000;
      20'h018d3: out <= 12'h000;
      20'h018d4: out <= 12'hfff;
      20'h018d5: out <= 12'h666;
      20'h018d6: out <= 12'h666;
      20'h018d7: out <= 12'h666;
      20'h018d8: out <= 12'h666;
      20'h018d9: out <= 12'h666;
      20'h018da: out <= 12'h666;
      20'h018db: out <= 12'h666;
      20'h018dc: out <= 12'hfff;
      20'h018dd: out <= 12'h666;
      20'h018de: out <= 12'h666;
      20'h018df: out <= 12'h666;
      20'h018e0: out <= 12'h666;
      20'h018e1: out <= 12'h666;
      20'h018e2: out <= 12'h666;
      20'h018e3: out <= 12'h666;
      20'h018e4: out <= 12'h603;
      20'h018e5: out <= 12'h603;
      20'h018e6: out <= 12'h603;
      20'h018e7: out <= 12'h603;
      20'h018e8: out <= 12'hee9;
      20'h018e9: out <= 12'hf87;
      20'h018ea: out <= 12'hf87;
      20'h018eb: out <= 12'hf87;
      20'h018ec: out <= 12'hf87;
      20'h018ed: out <= 12'hf87;
      20'h018ee: out <= 12'hf87;
      20'h018ef: out <= 12'hb27;
      20'h018f0: out <= 12'h000;
      20'h018f1: out <= 12'h000;
      20'h018f2: out <= 12'h000;
      20'h018f3: out <= 12'h000;
      20'h018f4: out <= 12'h000;
      20'h018f5: out <= 12'h000;
      20'h018f6: out <= 12'h000;
      20'h018f7: out <= 12'h000;
      20'h018f8: out <= 12'h000;
      20'h018f9: out <= 12'hee9;
      20'h018fa: out <= 12'hee9;
      20'h018fb: out <= 12'hee9;
      20'h018fc: out <= 12'hee9;
      20'h018fd: out <= 12'h000;
      20'h018fe: out <= 12'h000;
      20'h018ff: out <= 12'h000;
      20'h01900: out <= 12'h000;
      20'h01901: out <= 12'hee9;
      20'h01902: out <= 12'hee9;
      20'h01903: out <= 12'h000;
      20'h01904: out <= 12'h000;
      20'h01905: out <= 12'h000;
      20'h01906: out <= 12'hee9;
      20'h01907: out <= 12'hee9;
      20'h01908: out <= 12'h000;
      20'h01909: out <= 12'h000;
      20'h0190a: out <= 12'hee9;
      20'h0190b: out <= 12'hee9;
      20'h0190c: out <= 12'h000;
      20'h0190d: out <= 12'h000;
      20'h0190e: out <= 12'hee9;
      20'h0190f: out <= 12'hee9;
      20'h01910: out <= 12'hee9;
      20'h01911: out <= 12'hee9;
      20'h01912: out <= 12'h000;
      20'h01913: out <= 12'h000;
      20'h01914: out <= 12'hee9;
      20'h01915: out <= 12'hee9;
      20'h01916: out <= 12'hee9;
      20'h01917: out <= 12'hee9;
      20'h01918: out <= 12'hee9;
      20'h01919: out <= 12'h000;
      20'h0191a: out <= 12'h000;
      20'h0191b: out <= 12'h000;
      20'h0191c: out <= 12'h000;
      20'h0191d: out <= 12'h000;
      20'h0191e: out <= 12'h000;
      20'h0191f: out <= 12'h000;
      20'h01920: out <= 12'h000;
      20'h01921: out <= 12'h000;
      20'h01922: out <= 12'h000;
      20'h01923: out <= 12'h000;
      20'h01924: out <= 12'h000;
      20'h01925: out <= 12'h000;
      20'h01926: out <= 12'h000;
      20'h01927: out <= 12'h000;
      20'h01928: out <= 12'hfff;
      20'h01929: out <= 12'h6af;
      20'h0192a: out <= 12'h16d;
      20'h0192b: out <= 12'hfff;
      20'h0192c: out <= 12'h16d;
      20'h0192d: out <= 12'hfff;
      20'h0192e: out <= 12'hfff;
      20'h0192f: out <= 12'hfff;
      20'h01930: out <= 12'hfff;
      20'h01931: out <= 12'h16d;
      20'h01932: out <= 12'h16d;
      20'h01933: out <= 12'h6af;
      20'h01934: out <= 12'hfff;
      20'h01935: out <= 12'hfff;
      20'h01936: out <= 12'hfff;
      20'h01937: out <= 12'hfff;
      20'h01938: out <= 12'h16d;
      20'h01939: out <= 12'h6af;
      20'h0193a: out <= 12'hfff;
      20'h0193b: out <= 12'hfff;
      20'h0193c: out <= 12'h16d;
      20'h0193d: out <= 12'hfff;
      20'h0193e: out <= 12'hfff;
      20'h0193f: out <= 12'hfff;
      20'h01940: out <= 12'hfff;
      20'h01941: out <= 12'h16d;
      20'h01942: out <= 12'hfff;
      20'h01943: out <= 12'h6af;
      20'h01944: out <= 12'h16d;
      20'h01945: out <= 12'hfff;
      20'h01946: out <= 12'hfff;
      20'h01947: out <= 12'hfff;
      20'h01948: out <= 12'h000;
      20'h01949: out <= 12'hfff;
      20'h0194a: out <= 12'h6af;
      20'h0194b: out <= 12'h16d;
      20'h0194c: out <= 12'h16d;
      20'h0194d: out <= 12'h16d;
      20'h0194e: out <= 12'h16d;
      20'h0194f: out <= 12'h6af;
      20'h01950: out <= 12'hfff;
      20'h01951: out <= 12'h6af;
      20'h01952: out <= 12'h16d;
      20'h01953: out <= 12'h16d;
      20'h01954: out <= 12'h16d;
      20'h01955: out <= 12'h16d;
      20'h01956: out <= 12'h6af;
      20'h01957: out <= 12'hfff;
      20'h01958: out <= 12'h222;
      20'h01959: out <= 12'h16d;
      20'h0195a: out <= 12'h6af;
      20'h0195b: out <= 12'hfff;
      20'h0195c: out <= 12'h16d;
      20'h0195d: out <= 12'h16d;
      20'h0195e: out <= 12'h16d;
      20'h0195f: out <= 12'h6af;
      20'h01960: out <= 12'hfff;
      20'h01961: out <= 12'h6af;
      20'h01962: out <= 12'h16d;
      20'h01963: out <= 12'h16d;
      20'h01964: out <= 12'h16d;
      20'h01965: out <= 12'hfff;
      20'h01966: out <= 12'h6af;
      20'h01967: out <= 12'h16d;
      20'h01968: out <= 12'hfff;
      20'h01969: out <= 12'hfff;
      20'h0196a: out <= 12'hfff;
      20'h0196b: out <= 12'hfff;
      20'h0196c: out <= 12'h6af;
      20'h0196d: out <= 12'h16d;
      20'h0196e: out <= 12'h16d;
      20'h0196f: out <= 12'hfff;
      20'h01970: out <= 12'hfff;
      20'h01971: out <= 12'hfff;
      20'h01972: out <= 12'hfff;
      20'h01973: out <= 12'h16d;
      20'h01974: out <= 12'hfff;
      20'h01975: out <= 12'h16d;
      20'h01976: out <= 12'h6af;
      20'h01977: out <= 12'hfff;
      20'h01978: out <= 12'hfff;
      20'h01979: out <= 12'hfff;
      20'h0197a: out <= 12'hfff;
      20'h0197b: out <= 12'h16d;
      20'h0197c: out <= 12'h6af;
      20'h0197d: out <= 12'hfff;
      20'h0197e: out <= 12'h16d;
      20'h0197f: out <= 12'hfff;
      20'h01980: out <= 12'hfff;
      20'h01981: out <= 12'hfff;
      20'h01982: out <= 12'hfff;
      20'h01983: out <= 12'h16d;
      20'h01984: out <= 12'hfff;
      20'h01985: out <= 12'hfff;
      20'h01986: out <= 12'h6af;
      20'h01987: out <= 12'h16d;
      20'h01988: out <= 12'h000;
      20'h01989: out <= 12'hfff;
      20'h0198a: out <= 12'h6af;
      20'h0198b: out <= 12'h16d;
      20'h0198c: out <= 12'h16d;
      20'h0198d: out <= 12'h16d;
      20'h0198e: out <= 12'h6af;
      20'h0198f: out <= 12'hfff;
      20'h01990: out <= 12'hfff;
      20'h01991: out <= 12'hfff;
      20'h01992: out <= 12'h6af;
      20'h01993: out <= 12'h16d;
      20'h01994: out <= 12'h16d;
      20'h01995: out <= 12'h16d;
      20'h01996: out <= 12'h6af;
      20'h01997: out <= 12'hfff;
      20'h01998: out <= 12'h222;
      20'h01999: out <= 12'h16d;
      20'h0199a: out <= 12'h6af;
      20'h0199b: out <= 12'hfff;
      20'h0199c: out <= 12'h16d;
      20'h0199d: out <= 12'h16d;
      20'h0199e: out <= 12'h6af;
      20'h0199f: out <= 12'hfff;
      20'h019a0: out <= 12'hfff;
      20'h019a1: out <= 12'hfff;
      20'h019a2: out <= 12'h6af;
      20'h019a3: out <= 12'h16d;
      20'h019a4: out <= 12'h16d;
      20'h019a5: out <= 12'hfff;
      20'h019a6: out <= 12'h6af;
      20'h019a7: out <= 12'h16d;
      20'h019a8: out <= 12'h603;
      20'h019a9: out <= 12'h603;
      20'h019aa: out <= 12'h603;
      20'h019ab: out <= 12'h603;
      20'h019ac: out <= 12'h666;
      20'h019ad: out <= 12'h666;
      20'h019ae: out <= 12'h666;
      20'h019af: out <= 12'h666;
      20'h019b0: out <= 12'h666;
      20'h019b1: out <= 12'h666;
      20'h019b2: out <= 12'h666;
      20'h019b3: out <= 12'h666;
      20'h019b4: out <= 12'h666;
      20'h019b5: out <= 12'h666;
      20'h019b6: out <= 12'h666;
      20'h019b7: out <= 12'h666;
      20'h019b8: out <= 12'h666;
      20'h019b9: out <= 12'h666;
      20'h019ba: out <= 12'h666;
      20'h019bb: out <= 12'h666;
      20'h019bc: out <= 12'h000;
      20'h019bd: out <= 12'h000;
      20'h019be: out <= 12'h000;
      20'h019bf: out <= 12'h000;
      20'h019c0: out <= 12'h000;
      20'h019c1: out <= 12'h000;
      20'h019c2: out <= 12'h000;
      20'h019c3: out <= 12'h000;
      20'h019c4: out <= 12'h666;
      20'h019c5: out <= 12'h666;
      20'h019c6: out <= 12'h666;
      20'h019c7: out <= 12'h666;
      20'h019c8: out <= 12'h666;
      20'h019c9: out <= 12'h666;
      20'h019ca: out <= 12'h666;
      20'h019cb: out <= 12'h666;
      20'h019cc: out <= 12'h000;
      20'h019cd: out <= 12'h000;
      20'h019ce: out <= 12'h000;
      20'h019cf: out <= 12'h000;
      20'h019d0: out <= 12'h000;
      20'h019d1: out <= 12'h000;
      20'h019d2: out <= 12'h000;
      20'h019d3: out <= 12'h000;
      20'h019d4: out <= 12'h000;
      20'h019d5: out <= 12'h000;
      20'h019d6: out <= 12'h000;
      20'h019d7: out <= 12'h000;
      20'h019d8: out <= 12'h000;
      20'h019d9: out <= 12'h000;
      20'h019da: out <= 12'h000;
      20'h019db: out <= 12'h000;
      20'h019dc: out <= 12'h666;
      20'h019dd: out <= 12'h666;
      20'h019de: out <= 12'h666;
      20'h019df: out <= 12'h666;
      20'h019e0: out <= 12'h666;
      20'h019e1: out <= 12'h666;
      20'h019e2: out <= 12'h666;
      20'h019e3: out <= 12'h666;
      20'h019e4: out <= 12'h000;
      20'h019e5: out <= 12'h000;
      20'h019e6: out <= 12'h000;
      20'h019e7: out <= 12'h000;
      20'h019e8: out <= 12'h000;
      20'h019e9: out <= 12'h000;
      20'h019ea: out <= 12'h000;
      20'h019eb: out <= 12'h000;
      20'h019ec: out <= 12'h666;
      20'h019ed: out <= 12'h666;
      20'h019ee: out <= 12'h666;
      20'h019ef: out <= 12'h666;
      20'h019f0: out <= 12'h666;
      20'h019f1: out <= 12'h666;
      20'h019f2: out <= 12'h666;
      20'h019f3: out <= 12'h666;
      20'h019f4: out <= 12'h666;
      20'h019f5: out <= 12'h666;
      20'h019f6: out <= 12'h666;
      20'h019f7: out <= 12'h666;
      20'h019f8: out <= 12'h666;
      20'h019f9: out <= 12'h666;
      20'h019fa: out <= 12'h666;
      20'h019fb: out <= 12'h666;
      20'h019fc: out <= 12'h603;
      20'h019fd: out <= 12'h603;
      20'h019fe: out <= 12'h603;
      20'h019ff: out <= 12'h603;
      20'h01a00: out <= 12'hb27;
      20'h01a01: out <= 12'hb27;
      20'h01a02: out <= 12'hb27;
      20'h01a03: out <= 12'hb27;
      20'h01a04: out <= 12'hb27;
      20'h01a05: out <= 12'hb27;
      20'h01a06: out <= 12'hb27;
      20'h01a07: out <= 12'hb27;
      20'h01a08: out <= 12'h000;
      20'h01a09: out <= 12'h000;
      20'h01a0a: out <= 12'h000;
      20'h01a0b: out <= 12'h000;
      20'h01a0c: out <= 12'h000;
      20'h01a0d: out <= 12'h000;
      20'h01a0e: out <= 12'h000;
      20'h01a0f: out <= 12'h000;
      20'h01a10: out <= 12'h000;
      20'h01a11: out <= 12'h000;
      20'h01a12: out <= 12'h000;
      20'h01a13: out <= 12'h000;
      20'h01a14: out <= 12'h000;
      20'h01a15: out <= 12'h000;
      20'h01a16: out <= 12'h000;
      20'h01a17: out <= 12'h000;
      20'h01a18: out <= 12'h000;
      20'h01a19: out <= 12'h000;
      20'h01a1a: out <= 12'h000;
      20'h01a1b: out <= 12'h000;
      20'h01a1c: out <= 12'h000;
      20'h01a1d: out <= 12'h000;
      20'h01a1e: out <= 12'h000;
      20'h01a1f: out <= 12'h000;
      20'h01a20: out <= 12'h000;
      20'h01a21: out <= 12'h000;
      20'h01a22: out <= 12'h000;
      20'h01a23: out <= 12'h000;
      20'h01a24: out <= 12'h000;
      20'h01a25: out <= 12'h000;
      20'h01a26: out <= 12'h000;
      20'h01a27: out <= 12'h000;
      20'h01a28: out <= 12'h000;
      20'h01a29: out <= 12'h000;
      20'h01a2a: out <= 12'h000;
      20'h01a2b: out <= 12'h000;
      20'h01a2c: out <= 12'h000;
      20'h01a2d: out <= 12'h000;
      20'h01a2e: out <= 12'h000;
      20'h01a2f: out <= 12'h000;
      20'h01a30: out <= 12'h000;
      20'h01a31: out <= 12'h000;
      20'h01a32: out <= 12'h000;
      20'h01a33: out <= 12'h000;
      20'h01a34: out <= 12'h000;
      20'h01a35: out <= 12'h000;
      20'h01a36: out <= 12'h000;
      20'h01a37: out <= 12'h000;
      20'h01a38: out <= 12'h000;
      20'h01a39: out <= 12'h000;
      20'h01a3a: out <= 12'h000;
      20'h01a3b: out <= 12'h000;
      20'h01a3c: out <= 12'h000;
      20'h01a3d: out <= 12'h000;
      20'h01a3e: out <= 12'h000;
      20'h01a3f: out <= 12'h000;
      20'h01a40: out <= 12'hfff;
      20'h01a41: out <= 12'h6af;
      20'h01a42: out <= 12'h16d;
      20'h01a43: out <= 12'hfff;
      20'h01a44: out <= 12'h16d;
      20'h01a45: out <= 12'h6af;
      20'h01a46: out <= 12'hfff;
      20'h01a47: out <= 12'hfff;
      20'h01a48: out <= 12'h6af;
      20'h01a49: out <= 12'h16d;
      20'h01a4a: out <= 12'h16d;
      20'h01a4b: out <= 12'h6af;
      20'h01a4c: out <= 12'hfff;
      20'h01a4d: out <= 12'h16d;
      20'h01a4e: out <= 12'h16d;
      20'h01a4f: out <= 12'h6af;
      20'h01a50: out <= 12'h16d;
      20'h01a51: out <= 12'h6af;
      20'h01a52: out <= 12'hfff;
      20'h01a53: out <= 12'hfff;
      20'h01a54: out <= 12'h16d;
      20'h01a55: out <= 12'h6af;
      20'h01a56: out <= 12'hfff;
      20'h01a57: out <= 12'hfff;
      20'h01a58: out <= 12'h6af;
      20'h01a59: out <= 12'h16d;
      20'h01a5a: out <= 12'hfff;
      20'h01a5b: out <= 12'h6af;
      20'h01a5c: out <= 12'h16d;
      20'h01a5d: out <= 12'h16d;
      20'h01a5e: out <= 12'h16d;
      20'h01a5f: out <= 12'h6af;
      20'h01a60: out <= 12'h000;
      20'h01a61: out <= 12'hfff;
      20'h01a62: out <= 12'h6af;
      20'h01a63: out <= 12'h16d;
      20'h01a64: out <= 12'h16d;
      20'h01a65: out <= 12'h16d;
      20'h01a66: out <= 12'h6af;
      20'h01a67: out <= 12'hfff;
      20'h01a68: out <= 12'hfff;
      20'h01a69: out <= 12'hfff;
      20'h01a6a: out <= 12'h6af;
      20'h01a6b: out <= 12'h16d;
      20'h01a6c: out <= 12'h16d;
      20'h01a6d: out <= 12'h16d;
      20'h01a6e: out <= 12'h6af;
      20'h01a6f: out <= 12'hfff;
      20'h01a70: out <= 12'h222;
      20'h01a71: out <= 12'h16d;
      20'h01a72: out <= 12'h6af;
      20'h01a73: out <= 12'hfff;
      20'h01a74: out <= 12'h16d;
      20'h01a75: out <= 12'h16d;
      20'h01a76: out <= 12'h6af;
      20'h01a77: out <= 12'hfff;
      20'h01a78: out <= 12'hfff;
      20'h01a79: out <= 12'hfff;
      20'h01a7a: out <= 12'h6af;
      20'h01a7b: out <= 12'h16d;
      20'h01a7c: out <= 12'h16d;
      20'h01a7d: out <= 12'hfff;
      20'h01a7e: out <= 12'h6af;
      20'h01a7f: out <= 12'h16d;
      20'h01a80: out <= 12'h6af;
      20'h01a81: out <= 12'h16d;
      20'h01a82: out <= 12'h16d;
      20'h01a83: out <= 12'hfff;
      20'h01a84: out <= 12'h6af;
      20'h01a85: out <= 12'h16d;
      20'h01a86: out <= 12'h16d;
      20'h01a87: out <= 12'h6af;
      20'h01a88: out <= 12'hfff;
      20'h01a89: out <= 12'hfff;
      20'h01a8a: out <= 12'h6af;
      20'h01a8b: out <= 12'h16d;
      20'h01a8c: out <= 12'hfff;
      20'h01a8d: out <= 12'h16d;
      20'h01a8e: out <= 12'h6af;
      20'h01a8f: out <= 12'hfff;
      20'h01a90: out <= 12'h6af;
      20'h01a91: out <= 12'h16d;
      20'h01a92: out <= 12'h16d;
      20'h01a93: out <= 12'h16d;
      20'h01a94: out <= 12'h6af;
      20'h01a95: out <= 12'hfff;
      20'h01a96: out <= 12'h16d;
      20'h01a97: out <= 12'h6af;
      20'h01a98: out <= 12'hfff;
      20'h01a99: out <= 12'hfff;
      20'h01a9a: out <= 12'h6af;
      20'h01a9b: out <= 12'h16d;
      20'h01a9c: out <= 12'hfff;
      20'h01a9d: out <= 12'hfff;
      20'h01a9e: out <= 12'h6af;
      20'h01a9f: out <= 12'h16d;
      20'h01aa0: out <= 12'h000;
      20'h01aa1: out <= 12'hfff;
      20'h01aa2: out <= 12'h6af;
      20'h01aa3: out <= 12'h16d;
      20'h01aa4: out <= 12'h16d;
      20'h01aa5: out <= 12'h16d;
      20'h01aa6: out <= 12'h16d;
      20'h01aa7: out <= 12'h6af;
      20'h01aa8: out <= 12'hfff;
      20'h01aa9: out <= 12'h6af;
      20'h01aaa: out <= 12'h16d;
      20'h01aab: out <= 12'h16d;
      20'h01aac: out <= 12'h16d;
      20'h01aad: out <= 12'h16d;
      20'h01aae: out <= 12'h6af;
      20'h01aaf: out <= 12'hfff;
      20'h01ab0: out <= 12'h222;
      20'h01ab1: out <= 12'h16d;
      20'h01ab2: out <= 12'h6af;
      20'h01ab3: out <= 12'hfff;
      20'h01ab4: out <= 12'h16d;
      20'h01ab5: out <= 12'h16d;
      20'h01ab6: out <= 12'h16d;
      20'h01ab7: out <= 12'h6af;
      20'h01ab8: out <= 12'hfff;
      20'h01ab9: out <= 12'h6af;
      20'h01aba: out <= 12'h16d;
      20'h01abb: out <= 12'h16d;
      20'h01abc: out <= 12'h16d;
      20'h01abd: out <= 12'hfff;
      20'h01abe: out <= 12'h6af;
      20'h01abf: out <= 12'h16d;
      20'h01ac0: out <= 12'h603;
      20'h01ac1: out <= 12'h603;
      20'h01ac2: out <= 12'h603;
      20'h01ac3: out <= 12'h603;
      20'h01ac4: out <= 12'hfff;
      20'h01ac5: out <= 12'hfff;
      20'h01ac6: out <= 12'hfff;
      20'h01ac7: out <= 12'hfff;
      20'h01ac8: out <= 12'hfff;
      20'h01ac9: out <= 12'hfff;
      20'h01aca: out <= 12'hfff;
      20'h01acb: out <= 12'h666;
      20'h01acc: out <= 12'hfff;
      20'h01acd: out <= 12'hfff;
      20'h01ace: out <= 12'hfff;
      20'h01acf: out <= 12'hfff;
      20'h01ad0: out <= 12'hfff;
      20'h01ad1: out <= 12'hfff;
      20'h01ad2: out <= 12'hfff;
      20'h01ad3: out <= 12'h666;
      20'h01ad4: out <= 12'h000;
      20'h01ad5: out <= 12'h000;
      20'h01ad6: out <= 12'h000;
      20'h01ad7: out <= 12'h000;
      20'h01ad8: out <= 12'h000;
      20'h01ad9: out <= 12'h000;
      20'h01ada: out <= 12'h000;
      20'h01adb: out <= 12'h000;
      20'h01adc: out <= 12'hfff;
      20'h01add: out <= 12'hfff;
      20'h01ade: out <= 12'hfff;
      20'h01adf: out <= 12'hfff;
      20'h01ae0: out <= 12'hfff;
      20'h01ae1: out <= 12'hfff;
      20'h01ae2: out <= 12'hfff;
      20'h01ae3: out <= 12'h666;
      20'h01ae4: out <= 12'hfff;
      20'h01ae5: out <= 12'hfff;
      20'h01ae6: out <= 12'hfff;
      20'h01ae7: out <= 12'hfff;
      20'h01ae8: out <= 12'hfff;
      20'h01ae9: out <= 12'hfff;
      20'h01aea: out <= 12'hfff;
      20'h01aeb: out <= 12'h666;
      20'h01aec: out <= 12'hfff;
      20'h01aed: out <= 12'hfff;
      20'h01aee: out <= 12'hfff;
      20'h01aef: out <= 12'hfff;
      20'h01af0: out <= 12'hfff;
      20'h01af1: out <= 12'hfff;
      20'h01af2: out <= 12'hfff;
      20'h01af3: out <= 12'h666;
      20'h01af4: out <= 12'hfff;
      20'h01af5: out <= 12'hfff;
      20'h01af6: out <= 12'hfff;
      20'h01af7: out <= 12'hfff;
      20'h01af8: out <= 12'hfff;
      20'h01af9: out <= 12'hfff;
      20'h01afa: out <= 12'hfff;
      20'h01afb: out <= 12'h666;
      20'h01afc: out <= 12'h000;
      20'h01afd: out <= 12'h000;
      20'h01afe: out <= 12'h000;
      20'h01aff: out <= 12'h000;
      20'h01b00: out <= 12'h000;
      20'h01b01: out <= 12'h000;
      20'h01b02: out <= 12'h000;
      20'h01b03: out <= 12'h000;
      20'h01b04: out <= 12'h000;
      20'h01b05: out <= 12'h000;
      20'h01b06: out <= 12'h000;
      20'h01b07: out <= 12'h000;
      20'h01b08: out <= 12'h000;
      20'h01b09: out <= 12'h000;
      20'h01b0a: out <= 12'h000;
      20'h01b0b: out <= 12'h000;
      20'h01b0c: out <= 12'h000;
      20'h01b0d: out <= 12'h000;
      20'h01b0e: out <= 12'h000;
      20'h01b0f: out <= 12'h000;
      20'h01b10: out <= 12'h000;
      20'h01b11: out <= 12'h000;
      20'h01b12: out <= 12'h000;
      20'h01b13: out <= 12'h000;
      20'h01b14: out <= 12'h603;
      20'h01b15: out <= 12'h603;
      20'h01b16: out <= 12'h603;
      20'h01b17: out <= 12'h603;
      20'h01b18: out <= 12'hee9;
      20'h01b19: out <= 12'hee9;
      20'h01b1a: out <= 12'hee9;
      20'h01b1b: out <= 12'hee9;
      20'h01b1c: out <= 12'hee9;
      20'h01b1d: out <= 12'hee9;
      20'h01b1e: out <= 12'hee9;
      20'h01b1f: out <= 12'hb27;
      20'h01b20: out <= 12'h000;
      20'h01b21: out <= 12'h000;
      20'h01b22: out <= 12'h000;
      20'h01b23: out <= 12'h000;
      20'h01b24: out <= 12'h000;
      20'h01b25: out <= 12'h000;
      20'h01b26: out <= 12'h000;
      20'h01b27: out <= 12'h000;
      20'h01b28: out <= 12'h000;
      20'h01b29: out <= 12'h000;
      20'h01b2a: out <= 12'h000;
      20'h01b2b: out <= 12'h000;
      20'h01b2c: out <= 12'h000;
      20'h01b2d: out <= 12'h000;
      20'h01b2e: out <= 12'h000;
      20'h01b2f: out <= 12'h000;
      20'h01b30: out <= 12'h000;
      20'h01b31: out <= 12'h000;
      20'h01b32: out <= 12'h000;
      20'h01b33: out <= 12'h000;
      20'h01b34: out <= 12'h000;
      20'h01b35: out <= 12'h000;
      20'h01b36: out <= 12'h000;
      20'h01b37: out <= 12'h000;
      20'h01b38: out <= 12'h000;
      20'h01b39: out <= 12'h000;
      20'h01b3a: out <= 12'h000;
      20'h01b3b: out <= 12'h000;
      20'h01b3c: out <= 12'h000;
      20'h01b3d: out <= 12'h000;
      20'h01b3e: out <= 12'h000;
      20'h01b3f: out <= 12'h000;
      20'h01b40: out <= 12'h000;
      20'h01b41: out <= 12'h000;
      20'h01b42: out <= 12'h000;
      20'h01b43: out <= 12'h000;
      20'h01b44: out <= 12'h000;
      20'h01b45: out <= 12'h000;
      20'h01b46: out <= 12'h000;
      20'h01b47: out <= 12'h000;
      20'h01b48: out <= 12'h000;
      20'h01b49: out <= 12'h000;
      20'h01b4a: out <= 12'h000;
      20'h01b4b: out <= 12'h000;
      20'h01b4c: out <= 12'h000;
      20'h01b4d: out <= 12'h000;
      20'h01b4e: out <= 12'h000;
      20'h01b4f: out <= 12'h000;
      20'h01b50: out <= 12'h000;
      20'h01b51: out <= 12'h000;
      20'h01b52: out <= 12'h000;
      20'h01b53: out <= 12'h000;
      20'h01b54: out <= 12'h000;
      20'h01b55: out <= 12'h000;
      20'h01b56: out <= 12'h000;
      20'h01b57: out <= 12'h000;
      20'h01b58: out <= 12'hfff;
      20'h01b59: out <= 12'h6af;
      20'h01b5a: out <= 12'h16d;
      20'h01b5b: out <= 12'h6af;
      20'h01b5c: out <= 12'h16d;
      20'h01b5d: out <= 12'h16d;
      20'h01b5e: out <= 12'h6af;
      20'h01b5f: out <= 12'h6af;
      20'h01b60: out <= 12'h16d;
      20'h01b61: out <= 12'h16d;
      20'h01b62: out <= 12'h16d;
      20'h01b63: out <= 12'h6af;
      20'h01b64: out <= 12'hfff;
      20'h01b65: out <= 12'h000;
      20'h01b66: out <= 12'h000;
      20'h01b67: out <= 12'h000;
      20'h01b68: out <= 12'h16d;
      20'h01b69: out <= 12'h6af;
      20'h01b6a: out <= 12'hfff;
      20'h01b6b: out <= 12'h6af;
      20'h01b6c: out <= 12'h16d;
      20'h01b6d: out <= 12'h16d;
      20'h01b6e: out <= 12'h6af;
      20'h01b6f: out <= 12'h6af;
      20'h01b70: out <= 12'h16d;
      20'h01b71: out <= 12'h16d;
      20'h01b72: out <= 12'hfff;
      20'h01b73: out <= 12'h6af;
      20'h01b74: out <= 12'h16d;
      20'h01b75: out <= 12'h222;
      20'h01b76: out <= 12'h222;
      20'h01b77: out <= 12'h222;
      20'h01b78: out <= 12'h000;
      20'h01b79: out <= 12'hfff;
      20'h01b7a: out <= 12'h6af;
      20'h01b7b: out <= 12'h16d;
      20'h01b7c: out <= 12'h16d;
      20'h01b7d: out <= 12'h16d;
      20'h01b7e: out <= 12'h6af;
      20'h01b7f: out <= 12'hfff;
      20'h01b80: out <= 12'hfff;
      20'h01b81: out <= 12'hfff;
      20'h01b82: out <= 12'h6af;
      20'h01b83: out <= 12'h16d;
      20'h01b84: out <= 12'h16d;
      20'h01b85: out <= 12'h16d;
      20'h01b86: out <= 12'h6af;
      20'h01b87: out <= 12'hfff;
      20'h01b88: out <= 12'h222;
      20'h01b89: out <= 12'h16d;
      20'h01b8a: out <= 12'h6af;
      20'h01b8b: out <= 12'hfff;
      20'h01b8c: out <= 12'h16d;
      20'h01b8d: out <= 12'h16d;
      20'h01b8e: out <= 12'h6af;
      20'h01b8f: out <= 12'hfff;
      20'h01b90: out <= 12'hfff;
      20'h01b91: out <= 12'hfff;
      20'h01b92: out <= 12'h6af;
      20'h01b93: out <= 12'h16d;
      20'h01b94: out <= 12'h16d;
      20'h01b95: out <= 12'hfff;
      20'h01b96: out <= 12'h6af;
      20'h01b97: out <= 12'h16d;
      20'h01b98: out <= 12'h000;
      20'h01b99: out <= 12'h000;
      20'h01b9a: out <= 12'h000;
      20'h01b9b: out <= 12'hfff;
      20'h01b9c: out <= 12'h6af;
      20'h01b9d: out <= 12'h16d;
      20'h01b9e: out <= 12'h16d;
      20'h01b9f: out <= 12'h16d;
      20'h01ba0: out <= 12'h6af;
      20'h01ba1: out <= 12'h6af;
      20'h01ba2: out <= 12'h16d;
      20'h01ba3: out <= 12'h16d;
      20'h01ba4: out <= 12'h6af;
      20'h01ba5: out <= 12'h16d;
      20'h01ba6: out <= 12'h6af;
      20'h01ba7: out <= 12'hfff;
      20'h01ba8: out <= 12'h222;
      20'h01ba9: out <= 12'h222;
      20'h01baa: out <= 12'h222;
      20'h01bab: out <= 12'h16d;
      20'h01bac: out <= 12'h6af;
      20'h01bad: out <= 12'hfff;
      20'h01bae: out <= 12'h16d;
      20'h01baf: out <= 12'h16d;
      20'h01bb0: out <= 12'h6af;
      20'h01bb1: out <= 12'h6af;
      20'h01bb2: out <= 12'h16d;
      20'h01bb3: out <= 12'h16d;
      20'h01bb4: out <= 12'h6af;
      20'h01bb5: out <= 12'hfff;
      20'h01bb6: out <= 12'h6af;
      20'h01bb7: out <= 12'h16d;
      20'h01bb8: out <= 12'h000;
      20'h01bb9: out <= 12'h6af;
      20'h01bba: out <= 12'hfff;
      20'h01bbb: out <= 12'h6af;
      20'h01bbc: out <= 12'h16d;
      20'h01bbd: out <= 12'h16d;
      20'h01bbe: out <= 12'h16d;
      20'h01bbf: out <= 12'h16d;
      20'h01bc0: out <= 12'h16d;
      20'h01bc1: out <= 12'h16d;
      20'h01bc2: out <= 12'h16d;
      20'h01bc3: out <= 12'h16d;
      20'h01bc4: out <= 12'h16d;
      20'h01bc5: out <= 12'h6af;
      20'h01bc6: out <= 12'hfff;
      20'h01bc7: out <= 12'h6af;
      20'h01bc8: out <= 12'h222;
      20'h01bc9: out <= 12'h6af;
      20'h01bca: out <= 12'h16d;
      20'h01bcb: out <= 12'h6af;
      20'h01bcc: out <= 12'hfff;
      20'h01bcd: out <= 12'hfff;
      20'h01bce: out <= 12'h16d;
      20'h01bcf: out <= 12'h16d;
      20'h01bd0: out <= 12'h16d;
      20'h01bd1: out <= 12'h16d;
      20'h01bd2: out <= 12'h16d;
      20'h01bd3: out <= 12'hfff;
      20'h01bd4: out <= 12'hfff;
      20'h01bd5: out <= 12'h6af;
      20'h01bd6: out <= 12'h16d;
      20'h01bd7: out <= 12'h6af;
      20'h01bd8: out <= 12'h603;
      20'h01bd9: out <= 12'h603;
      20'h01bda: out <= 12'h603;
      20'h01bdb: out <= 12'h603;
      20'h01bdc: out <= 12'hfff;
      20'h01bdd: out <= 12'hbbb;
      20'h01bde: out <= 12'hbbb;
      20'h01bdf: out <= 12'hbbb;
      20'h01be0: out <= 12'hbbb;
      20'h01be1: out <= 12'hbbb;
      20'h01be2: out <= 12'h666;
      20'h01be3: out <= 12'h666;
      20'h01be4: out <= 12'hfff;
      20'h01be5: out <= 12'hbbb;
      20'h01be6: out <= 12'hbbb;
      20'h01be7: out <= 12'hbbb;
      20'h01be8: out <= 12'hbbb;
      20'h01be9: out <= 12'hbbb;
      20'h01bea: out <= 12'h666;
      20'h01beb: out <= 12'h666;
      20'h01bec: out <= 12'h000;
      20'h01bed: out <= 12'h000;
      20'h01bee: out <= 12'h000;
      20'h01bef: out <= 12'h000;
      20'h01bf0: out <= 12'h000;
      20'h01bf1: out <= 12'h000;
      20'h01bf2: out <= 12'h000;
      20'h01bf3: out <= 12'h000;
      20'h01bf4: out <= 12'hfff;
      20'h01bf5: out <= 12'hbbb;
      20'h01bf6: out <= 12'hbbb;
      20'h01bf7: out <= 12'hbbb;
      20'h01bf8: out <= 12'hbbb;
      20'h01bf9: out <= 12'hbbb;
      20'h01bfa: out <= 12'h666;
      20'h01bfb: out <= 12'h666;
      20'h01bfc: out <= 12'hfff;
      20'h01bfd: out <= 12'hbbb;
      20'h01bfe: out <= 12'hbbb;
      20'h01bff: out <= 12'hbbb;
      20'h01c00: out <= 12'hbbb;
      20'h01c01: out <= 12'hbbb;
      20'h01c02: out <= 12'h666;
      20'h01c03: out <= 12'h666;
      20'h01c04: out <= 12'hfff;
      20'h01c05: out <= 12'hbbb;
      20'h01c06: out <= 12'hbbb;
      20'h01c07: out <= 12'hbbb;
      20'h01c08: out <= 12'hbbb;
      20'h01c09: out <= 12'hbbb;
      20'h01c0a: out <= 12'h666;
      20'h01c0b: out <= 12'h666;
      20'h01c0c: out <= 12'hfff;
      20'h01c0d: out <= 12'hbbb;
      20'h01c0e: out <= 12'hbbb;
      20'h01c0f: out <= 12'hbbb;
      20'h01c10: out <= 12'hbbb;
      20'h01c11: out <= 12'hbbb;
      20'h01c12: out <= 12'h666;
      20'h01c13: out <= 12'h666;
      20'h01c14: out <= 12'h000;
      20'h01c15: out <= 12'h000;
      20'h01c16: out <= 12'h000;
      20'h01c17: out <= 12'h000;
      20'h01c18: out <= 12'h000;
      20'h01c19: out <= 12'h000;
      20'h01c1a: out <= 12'h000;
      20'h01c1b: out <= 12'h000;
      20'h01c1c: out <= 12'h000;
      20'h01c1d: out <= 12'h000;
      20'h01c1e: out <= 12'h000;
      20'h01c1f: out <= 12'h000;
      20'h01c20: out <= 12'h000;
      20'h01c21: out <= 12'h000;
      20'h01c22: out <= 12'h000;
      20'h01c23: out <= 12'h000;
      20'h01c24: out <= 12'h000;
      20'h01c25: out <= 12'h000;
      20'h01c26: out <= 12'h000;
      20'h01c27: out <= 12'h000;
      20'h01c28: out <= 12'h000;
      20'h01c29: out <= 12'h000;
      20'h01c2a: out <= 12'h000;
      20'h01c2b: out <= 12'h000;
      20'h01c2c: out <= 12'h603;
      20'h01c2d: out <= 12'h603;
      20'h01c2e: out <= 12'h603;
      20'h01c2f: out <= 12'h603;
      20'h01c30: out <= 12'hee9;
      20'h01c31: out <= 12'hf87;
      20'h01c32: out <= 12'hf87;
      20'h01c33: out <= 12'hf87;
      20'h01c34: out <= 12'hf87;
      20'h01c35: out <= 12'hf87;
      20'h01c36: out <= 12'hf87;
      20'h01c37: out <= 12'hb27;
      20'h01c38: out <= 12'h000;
      20'h01c39: out <= 12'h000;
      20'h01c3a: out <= 12'h000;
      20'h01c3b: out <= 12'h000;
      20'h01c3c: out <= 12'h000;
      20'h01c3d: out <= 12'h000;
      20'h01c3e: out <= 12'h000;
      20'h01c3f: out <= 12'h000;
      20'h01c40: out <= 12'h000;
      20'h01c41: out <= 12'h000;
      20'h01c42: out <= 12'h000;
      20'h01c43: out <= 12'h000;
      20'h01c44: out <= 12'h000;
      20'h01c45: out <= 12'h000;
      20'h01c46: out <= 12'h000;
      20'h01c47: out <= 12'h000;
      20'h01c48: out <= 12'h000;
      20'h01c49: out <= 12'h000;
      20'h01c4a: out <= 12'h000;
      20'h01c4b: out <= 12'h000;
      20'h01c4c: out <= 12'h000;
      20'h01c4d: out <= 12'h000;
      20'h01c4e: out <= 12'h000;
      20'h01c4f: out <= 12'h000;
      20'h01c50: out <= 12'h000;
      20'h01c51: out <= 12'h000;
      20'h01c52: out <= 12'h000;
      20'h01c53: out <= 12'h000;
      20'h01c54: out <= 12'h000;
      20'h01c55: out <= 12'h000;
      20'h01c56: out <= 12'h000;
      20'h01c57: out <= 12'h000;
      20'h01c58: out <= 12'h000;
      20'h01c59: out <= 12'h000;
      20'h01c5a: out <= 12'h000;
      20'h01c5b: out <= 12'h000;
      20'h01c5c: out <= 12'h000;
      20'h01c5d: out <= 12'h000;
      20'h01c5e: out <= 12'h000;
      20'h01c5f: out <= 12'h000;
      20'h01c60: out <= 12'h000;
      20'h01c61: out <= 12'h000;
      20'h01c62: out <= 12'h000;
      20'h01c63: out <= 12'h000;
      20'h01c64: out <= 12'h000;
      20'h01c65: out <= 12'h000;
      20'h01c66: out <= 12'h000;
      20'h01c67: out <= 12'h000;
      20'h01c68: out <= 12'h000;
      20'h01c69: out <= 12'h000;
      20'h01c6a: out <= 12'h000;
      20'h01c6b: out <= 12'h000;
      20'h01c6c: out <= 12'h000;
      20'h01c6d: out <= 12'h000;
      20'h01c6e: out <= 12'h000;
      20'h01c6f: out <= 12'h000;
      20'h01c70: out <= 12'h000;
      20'h01c71: out <= 12'hfff;
      20'h01c72: out <= 12'h6af;
      20'h01c73: out <= 12'h16d;
      20'h01c74: out <= 12'h6af;
      20'h01c75: out <= 12'h16d;
      20'h01c76: out <= 12'h16d;
      20'h01c77: out <= 12'h16d;
      20'h01c78: out <= 12'h16d;
      20'h01c79: out <= 12'h16d;
      20'h01c7a: out <= 12'h6af;
      20'h01c7b: out <= 12'hfff;
      20'h01c7c: out <= 12'h000;
      20'h01c7d: out <= 12'h000;
      20'h01c7e: out <= 12'h000;
      20'h01c7f: out <= 12'h000;
      20'h01c80: out <= 12'h222;
      20'h01c81: out <= 12'h16d;
      20'h01c82: out <= 12'h6af;
      20'h01c83: out <= 12'hfff;
      20'h01c84: out <= 12'h6af;
      20'h01c85: out <= 12'h16d;
      20'h01c86: out <= 12'h16d;
      20'h01c87: out <= 12'h16d;
      20'h01c88: out <= 12'h16d;
      20'h01c89: out <= 12'hfff;
      20'h01c8a: out <= 12'h6af;
      20'h01c8b: out <= 12'h16d;
      20'h01c8c: out <= 12'h222;
      20'h01c8d: out <= 12'h222;
      20'h01c8e: out <= 12'h222;
      20'h01c8f: out <= 12'h222;
      20'h01c90: out <= 12'h000;
      20'h01c91: out <= 12'hfff;
      20'h01c92: out <= 12'h6af;
      20'h01c93: out <= 12'h16d;
      20'h01c94: out <= 12'h16d;
      20'h01c95: out <= 12'h16d;
      20'h01c96: out <= 12'h16d;
      20'h01c97: out <= 12'h6af;
      20'h01c98: out <= 12'hfff;
      20'h01c99: out <= 12'h6af;
      20'h01c9a: out <= 12'h16d;
      20'h01c9b: out <= 12'h16d;
      20'h01c9c: out <= 12'h16d;
      20'h01c9d: out <= 12'h16d;
      20'h01c9e: out <= 12'h6af;
      20'h01c9f: out <= 12'hfff;
      20'h01ca0: out <= 12'h222;
      20'h01ca1: out <= 12'h16d;
      20'h01ca2: out <= 12'h6af;
      20'h01ca3: out <= 12'hfff;
      20'h01ca4: out <= 12'h16d;
      20'h01ca5: out <= 12'h16d;
      20'h01ca6: out <= 12'h16d;
      20'h01ca7: out <= 12'h6af;
      20'h01ca8: out <= 12'hfff;
      20'h01ca9: out <= 12'h6af;
      20'h01caa: out <= 12'h16d;
      20'h01cab: out <= 12'h16d;
      20'h01cac: out <= 12'h16d;
      20'h01cad: out <= 12'hfff;
      20'h01cae: out <= 12'h6af;
      20'h01caf: out <= 12'h16d;
      20'h01cb0: out <= 12'h000;
      20'h01cb1: out <= 12'h000;
      20'h01cb2: out <= 12'h000;
      20'h01cb3: out <= 12'h000;
      20'h01cb4: out <= 12'hfff;
      20'h01cb5: out <= 12'h6af;
      20'h01cb6: out <= 12'h16d;
      20'h01cb7: out <= 12'h16d;
      20'h01cb8: out <= 12'h16d;
      20'h01cb9: out <= 12'h16d;
      20'h01cba: out <= 12'h16d;
      20'h01cbb: out <= 12'h6af;
      20'h01cbc: out <= 12'h16d;
      20'h01cbd: out <= 12'h6af;
      20'h01cbe: out <= 12'hfff;
      20'h01cbf: out <= 12'h000;
      20'h01cc0: out <= 12'h222;
      20'h01cc1: out <= 12'h222;
      20'h01cc2: out <= 12'h222;
      20'h01cc3: out <= 12'h222;
      20'h01cc4: out <= 12'h16d;
      20'h01cc5: out <= 12'h6af;
      20'h01cc6: out <= 12'hfff;
      20'h01cc7: out <= 12'h16d;
      20'h01cc8: out <= 12'h16d;
      20'h01cc9: out <= 12'h16d;
      20'h01cca: out <= 12'h16d;
      20'h01ccb: out <= 12'h6af;
      20'h01ccc: out <= 12'hfff;
      20'h01ccd: out <= 12'h6af;
      20'h01cce: out <= 12'h16d;
      20'h01ccf: out <= 12'h222;
      20'h01cd0: out <= 12'h000;
      20'h01cd1: out <= 12'h6af;
      20'h01cd2: out <= 12'h16d;
      20'h01cd3: out <= 12'hfff;
      20'h01cd4: out <= 12'h6af;
      20'h01cd5: out <= 12'h6af;
      20'h01cd6: out <= 12'h16d;
      20'h01cd7: out <= 12'h16d;
      20'h01cd8: out <= 12'h16d;
      20'h01cd9: out <= 12'h16d;
      20'h01cda: out <= 12'h16d;
      20'h01cdb: out <= 12'h6af;
      20'h01cdc: out <= 12'h6af;
      20'h01cdd: out <= 12'hfff;
      20'h01cde: out <= 12'h16d;
      20'h01cdf: out <= 12'h6af;
      20'h01ce0: out <= 12'h222;
      20'h01ce1: out <= 12'h6af;
      20'h01ce2: out <= 12'h16d;
      20'h01ce3: out <= 12'h16d;
      20'h01ce4: out <= 12'h6af;
      20'h01ce5: out <= 12'h6af;
      20'h01ce6: out <= 12'hfff;
      20'h01ce7: out <= 12'hfff;
      20'h01ce8: out <= 12'hfff;
      20'h01ce9: out <= 12'hfff;
      20'h01cea: out <= 12'hfff;
      20'h01ceb: out <= 12'h6af;
      20'h01cec: out <= 12'h6af;
      20'h01ced: out <= 12'h16d;
      20'h01cee: out <= 12'h16d;
      20'h01cef: out <= 12'h6af;
      20'h01cf0: out <= 12'h603;
      20'h01cf1: out <= 12'h603;
      20'h01cf2: out <= 12'h603;
      20'h01cf3: out <= 12'h603;
      20'h01cf4: out <= 12'hfff;
      20'h01cf5: out <= 12'hbbb;
      20'h01cf6: out <= 12'h666;
      20'h01cf7: out <= 12'h666;
      20'h01cf8: out <= 12'h666;
      20'h01cf9: out <= 12'hbbb;
      20'h01cfa: out <= 12'h666;
      20'h01cfb: out <= 12'h666;
      20'h01cfc: out <= 12'hfff;
      20'h01cfd: out <= 12'hbbb;
      20'h01cfe: out <= 12'h666;
      20'h01cff: out <= 12'h666;
      20'h01d00: out <= 12'h666;
      20'h01d01: out <= 12'hbbb;
      20'h01d02: out <= 12'h666;
      20'h01d03: out <= 12'h666;
      20'h01d04: out <= 12'h000;
      20'h01d05: out <= 12'h000;
      20'h01d06: out <= 12'h000;
      20'h01d07: out <= 12'h000;
      20'h01d08: out <= 12'h000;
      20'h01d09: out <= 12'h000;
      20'h01d0a: out <= 12'h000;
      20'h01d0b: out <= 12'h000;
      20'h01d0c: out <= 12'hfff;
      20'h01d0d: out <= 12'hbbb;
      20'h01d0e: out <= 12'h666;
      20'h01d0f: out <= 12'h666;
      20'h01d10: out <= 12'h666;
      20'h01d11: out <= 12'hbbb;
      20'h01d12: out <= 12'h666;
      20'h01d13: out <= 12'h666;
      20'h01d14: out <= 12'hfff;
      20'h01d15: out <= 12'hbbb;
      20'h01d16: out <= 12'h666;
      20'h01d17: out <= 12'h666;
      20'h01d18: out <= 12'h666;
      20'h01d19: out <= 12'hbbb;
      20'h01d1a: out <= 12'h666;
      20'h01d1b: out <= 12'h666;
      20'h01d1c: out <= 12'hfff;
      20'h01d1d: out <= 12'hbbb;
      20'h01d1e: out <= 12'h666;
      20'h01d1f: out <= 12'h666;
      20'h01d20: out <= 12'h666;
      20'h01d21: out <= 12'hbbb;
      20'h01d22: out <= 12'h666;
      20'h01d23: out <= 12'h666;
      20'h01d24: out <= 12'hfff;
      20'h01d25: out <= 12'hbbb;
      20'h01d26: out <= 12'h666;
      20'h01d27: out <= 12'h666;
      20'h01d28: out <= 12'h666;
      20'h01d29: out <= 12'hbbb;
      20'h01d2a: out <= 12'h666;
      20'h01d2b: out <= 12'h666;
      20'h01d2c: out <= 12'h000;
      20'h01d2d: out <= 12'h000;
      20'h01d2e: out <= 12'h000;
      20'h01d2f: out <= 12'h000;
      20'h01d30: out <= 12'h000;
      20'h01d31: out <= 12'h000;
      20'h01d32: out <= 12'h000;
      20'h01d33: out <= 12'h000;
      20'h01d34: out <= 12'h000;
      20'h01d35: out <= 12'h000;
      20'h01d36: out <= 12'h000;
      20'h01d37: out <= 12'h000;
      20'h01d38: out <= 12'h000;
      20'h01d39: out <= 12'h000;
      20'h01d3a: out <= 12'h000;
      20'h01d3b: out <= 12'h000;
      20'h01d3c: out <= 12'h000;
      20'h01d3d: out <= 12'h000;
      20'h01d3e: out <= 12'h000;
      20'h01d3f: out <= 12'h000;
      20'h01d40: out <= 12'h000;
      20'h01d41: out <= 12'h000;
      20'h01d42: out <= 12'h000;
      20'h01d43: out <= 12'h000;
      20'h01d44: out <= 12'h603;
      20'h01d45: out <= 12'h603;
      20'h01d46: out <= 12'h603;
      20'h01d47: out <= 12'h603;
      20'h01d48: out <= 12'hee9;
      20'h01d49: out <= 12'hf87;
      20'h01d4a: out <= 12'hee9;
      20'h01d4b: out <= 12'hee9;
      20'h01d4c: out <= 12'hee9;
      20'h01d4d: out <= 12'hb27;
      20'h01d4e: out <= 12'hf87;
      20'h01d4f: out <= 12'hb27;
      20'h01d50: out <= 12'h000;
      20'h01d51: out <= 12'h000;
      20'h01d52: out <= 12'h000;
      20'h01d53: out <= 12'h000;
      20'h01d54: out <= 12'h000;
      20'h01d55: out <= 12'h000;
      20'h01d56: out <= 12'h000;
      20'h01d57: out <= 12'h000;
      20'h01d58: out <= 12'h000;
      20'h01d59: out <= 12'h000;
      20'h01d5a: out <= 12'h000;
      20'h01d5b: out <= 12'h000;
      20'h01d5c: out <= 12'h000;
      20'h01d5d: out <= 12'h000;
      20'h01d5e: out <= 12'h000;
      20'h01d5f: out <= 12'h000;
      20'h01d60: out <= 12'h000;
      20'h01d61: out <= 12'h000;
      20'h01d62: out <= 12'h000;
      20'h01d63: out <= 12'h000;
      20'h01d64: out <= 12'h000;
      20'h01d65: out <= 12'h000;
      20'h01d66: out <= 12'h000;
      20'h01d67: out <= 12'h000;
      20'h01d68: out <= 12'h000;
      20'h01d69: out <= 12'h000;
      20'h01d6a: out <= 12'h000;
      20'h01d6b: out <= 12'h000;
      20'h01d6c: out <= 12'h000;
      20'h01d6d: out <= 12'h000;
      20'h01d6e: out <= 12'h000;
      20'h01d6f: out <= 12'h000;
      20'h01d70: out <= 12'h000;
      20'h01d71: out <= 12'h000;
      20'h01d72: out <= 12'h000;
      20'h01d73: out <= 12'h000;
      20'h01d74: out <= 12'h000;
      20'h01d75: out <= 12'h000;
      20'h01d76: out <= 12'h000;
      20'h01d77: out <= 12'h000;
      20'h01d78: out <= 12'h000;
      20'h01d79: out <= 12'h000;
      20'h01d7a: out <= 12'h000;
      20'h01d7b: out <= 12'h000;
      20'h01d7c: out <= 12'h000;
      20'h01d7d: out <= 12'h000;
      20'h01d7e: out <= 12'h000;
      20'h01d7f: out <= 12'h000;
      20'h01d80: out <= 12'h000;
      20'h01d81: out <= 12'h000;
      20'h01d82: out <= 12'h000;
      20'h01d83: out <= 12'h000;
      20'h01d84: out <= 12'h000;
      20'h01d85: out <= 12'h000;
      20'h01d86: out <= 12'h000;
      20'h01d87: out <= 12'h000;
      20'h01d88: out <= 12'h000;
      20'h01d89: out <= 12'hfff;
      20'h01d8a: out <= 12'h6af;
      20'h01d8b: out <= 12'h16d;
      20'h01d8c: out <= 12'h16d;
      20'h01d8d: out <= 12'h16d;
      20'h01d8e: out <= 12'h16d;
      20'h01d8f: out <= 12'h16d;
      20'h01d90: out <= 12'h16d;
      20'h01d91: out <= 12'h16d;
      20'h01d92: out <= 12'h6af;
      20'h01d93: out <= 12'hfff;
      20'h01d94: out <= 12'h000;
      20'h01d95: out <= 12'h000;
      20'h01d96: out <= 12'h000;
      20'h01d97: out <= 12'h000;
      20'h01d98: out <= 12'h222;
      20'h01d99: out <= 12'h16d;
      20'h01d9a: out <= 12'h6af;
      20'h01d9b: out <= 12'hfff;
      20'h01d9c: out <= 12'h16d;
      20'h01d9d: out <= 12'h16d;
      20'h01d9e: out <= 12'h16d;
      20'h01d9f: out <= 12'h16d;
      20'h01da0: out <= 12'h16d;
      20'h01da1: out <= 12'hfff;
      20'h01da2: out <= 12'h6af;
      20'h01da3: out <= 12'h16d;
      20'h01da4: out <= 12'h222;
      20'h01da5: out <= 12'h222;
      20'h01da6: out <= 12'h222;
      20'h01da7: out <= 12'h222;
      20'h01da8: out <= 12'h000;
      20'h01da9: out <= 12'hfff;
      20'h01daa: out <= 12'h6af;
      20'h01dab: out <= 12'h16d;
      20'h01dac: out <= 12'h16d;
      20'h01dad: out <= 12'h6af;
      20'h01dae: out <= 12'h16d;
      20'h01daf: out <= 12'h16d;
      20'h01db0: out <= 12'h16d;
      20'h01db1: out <= 12'h16d;
      20'h01db2: out <= 12'h16d;
      20'h01db3: out <= 12'h6af;
      20'h01db4: out <= 12'h16d;
      20'h01db5: out <= 12'h16d;
      20'h01db6: out <= 12'h6af;
      20'h01db7: out <= 12'hfff;
      20'h01db8: out <= 12'h222;
      20'h01db9: out <= 12'h16d;
      20'h01dba: out <= 12'h6af;
      20'h01dbb: out <= 12'hfff;
      20'h01dbc: out <= 12'h16d;
      20'h01dbd: out <= 12'h6af;
      20'h01dbe: out <= 12'h16d;
      20'h01dbf: out <= 12'h16d;
      20'h01dc0: out <= 12'h16d;
      20'h01dc1: out <= 12'h16d;
      20'h01dc2: out <= 12'h16d;
      20'h01dc3: out <= 12'h6af;
      20'h01dc4: out <= 12'h16d;
      20'h01dc5: out <= 12'hfff;
      20'h01dc6: out <= 12'h6af;
      20'h01dc7: out <= 12'h16d;
      20'h01dc8: out <= 12'h000;
      20'h01dc9: out <= 12'h000;
      20'h01dca: out <= 12'h000;
      20'h01dcb: out <= 12'h000;
      20'h01dcc: out <= 12'hfff;
      20'h01dcd: out <= 12'h6af;
      20'h01dce: out <= 12'h16d;
      20'h01dcf: out <= 12'h16d;
      20'h01dd0: out <= 12'h16d;
      20'h01dd1: out <= 12'h16d;
      20'h01dd2: out <= 12'h16d;
      20'h01dd3: out <= 12'h16d;
      20'h01dd4: out <= 12'h16d;
      20'h01dd5: out <= 12'h6af;
      20'h01dd6: out <= 12'hfff;
      20'h01dd7: out <= 12'h000;
      20'h01dd8: out <= 12'h222;
      20'h01dd9: out <= 12'h222;
      20'h01dda: out <= 12'h222;
      20'h01ddb: out <= 12'h222;
      20'h01ddc: out <= 12'h16d;
      20'h01ddd: out <= 12'h6af;
      20'h01dde: out <= 12'hfff;
      20'h01ddf: out <= 12'h16d;
      20'h01de0: out <= 12'h16d;
      20'h01de1: out <= 12'h16d;
      20'h01de2: out <= 12'h16d;
      20'h01de3: out <= 12'h16d;
      20'h01de4: out <= 12'hfff;
      20'h01de5: out <= 12'h6af;
      20'h01de6: out <= 12'h16d;
      20'h01de7: out <= 12'h222;
      20'h01de8: out <= 12'h000;
      20'h01de9: out <= 12'hfff;
      20'h01dea: out <= 12'hfff;
      20'h01deb: out <= 12'hfff;
      20'h01dec: out <= 12'hfff;
      20'h01ded: out <= 12'hfff;
      20'h01dee: out <= 12'h6af;
      20'h01def: out <= 12'h6af;
      20'h01df0: out <= 12'h6af;
      20'h01df1: out <= 12'h6af;
      20'h01df2: out <= 12'h6af;
      20'h01df3: out <= 12'hfff;
      20'h01df4: out <= 12'hfff;
      20'h01df5: out <= 12'hfff;
      20'h01df6: out <= 12'hfff;
      20'h01df7: out <= 12'hfff;
      20'h01df8: out <= 12'h222;
      20'h01df9: out <= 12'hfff;
      20'h01dfa: out <= 12'hfff;
      20'h01dfb: out <= 12'hfff;
      20'h01dfc: out <= 12'h16d;
      20'h01dfd: out <= 12'h16d;
      20'h01dfe: out <= 12'h6af;
      20'h01dff: out <= 12'h6af;
      20'h01e00: out <= 12'h6af;
      20'h01e01: out <= 12'h6af;
      20'h01e02: out <= 12'h6af;
      20'h01e03: out <= 12'h16d;
      20'h01e04: out <= 12'h16d;
      20'h01e05: out <= 12'hfff;
      20'h01e06: out <= 12'hfff;
      20'h01e07: out <= 12'hfff;
      20'h01e08: out <= 12'h603;
      20'h01e09: out <= 12'h603;
      20'h01e0a: out <= 12'h603;
      20'h01e0b: out <= 12'h603;
      20'h01e0c: out <= 12'hfff;
      20'h01e0d: out <= 12'hbbb;
      20'h01e0e: out <= 12'h666;
      20'h01e0f: out <= 12'hbbb;
      20'h01e10: out <= 12'hfff;
      20'h01e11: out <= 12'hbbb;
      20'h01e12: out <= 12'h666;
      20'h01e13: out <= 12'h666;
      20'h01e14: out <= 12'hfff;
      20'h01e15: out <= 12'hbbb;
      20'h01e16: out <= 12'h666;
      20'h01e17: out <= 12'hbbb;
      20'h01e18: out <= 12'hfff;
      20'h01e19: out <= 12'hbbb;
      20'h01e1a: out <= 12'h666;
      20'h01e1b: out <= 12'h666;
      20'h01e1c: out <= 12'h000;
      20'h01e1d: out <= 12'h000;
      20'h01e1e: out <= 12'h000;
      20'h01e1f: out <= 12'h000;
      20'h01e20: out <= 12'h000;
      20'h01e21: out <= 12'h000;
      20'h01e22: out <= 12'h000;
      20'h01e23: out <= 12'h000;
      20'h01e24: out <= 12'hfff;
      20'h01e25: out <= 12'hbbb;
      20'h01e26: out <= 12'h666;
      20'h01e27: out <= 12'hbbb;
      20'h01e28: out <= 12'hfff;
      20'h01e29: out <= 12'hbbb;
      20'h01e2a: out <= 12'h666;
      20'h01e2b: out <= 12'h666;
      20'h01e2c: out <= 12'hfff;
      20'h01e2d: out <= 12'hbbb;
      20'h01e2e: out <= 12'h666;
      20'h01e2f: out <= 12'hbbb;
      20'h01e30: out <= 12'hfff;
      20'h01e31: out <= 12'hbbb;
      20'h01e32: out <= 12'h666;
      20'h01e33: out <= 12'h666;
      20'h01e34: out <= 12'hfff;
      20'h01e35: out <= 12'hbbb;
      20'h01e36: out <= 12'h666;
      20'h01e37: out <= 12'hbbb;
      20'h01e38: out <= 12'hfff;
      20'h01e39: out <= 12'hbbb;
      20'h01e3a: out <= 12'h666;
      20'h01e3b: out <= 12'h666;
      20'h01e3c: out <= 12'hfff;
      20'h01e3d: out <= 12'hbbb;
      20'h01e3e: out <= 12'h666;
      20'h01e3f: out <= 12'hbbb;
      20'h01e40: out <= 12'hfff;
      20'h01e41: out <= 12'hbbb;
      20'h01e42: out <= 12'h666;
      20'h01e43: out <= 12'h666;
      20'h01e44: out <= 12'h000;
      20'h01e45: out <= 12'h000;
      20'h01e46: out <= 12'h000;
      20'h01e47: out <= 12'h000;
      20'h01e48: out <= 12'h000;
      20'h01e49: out <= 12'h000;
      20'h01e4a: out <= 12'h000;
      20'h01e4b: out <= 12'h000;
      20'h01e4c: out <= 12'h000;
      20'h01e4d: out <= 12'h000;
      20'h01e4e: out <= 12'h000;
      20'h01e4f: out <= 12'h000;
      20'h01e50: out <= 12'h000;
      20'h01e51: out <= 12'h000;
      20'h01e52: out <= 12'h000;
      20'h01e53: out <= 12'h000;
      20'h01e54: out <= 12'h000;
      20'h01e55: out <= 12'h000;
      20'h01e56: out <= 12'h000;
      20'h01e57: out <= 12'h000;
      20'h01e58: out <= 12'h000;
      20'h01e59: out <= 12'h000;
      20'h01e5a: out <= 12'h000;
      20'h01e5b: out <= 12'h000;
      20'h01e5c: out <= 12'h603;
      20'h01e5d: out <= 12'h603;
      20'h01e5e: out <= 12'h603;
      20'h01e5f: out <= 12'h603;
      20'h01e60: out <= 12'hee9;
      20'h01e61: out <= 12'hf87;
      20'h01e62: out <= 12'hee9;
      20'h01e63: out <= 12'hf87;
      20'h01e64: out <= 12'hf87;
      20'h01e65: out <= 12'hb27;
      20'h01e66: out <= 12'hf87;
      20'h01e67: out <= 12'hb27;
      20'h01e68: out <= 12'h000;
      20'h01e69: out <= 12'h000;
      20'h01e6a: out <= 12'h000;
      20'h01e6b: out <= 12'h000;
      20'h01e6c: out <= 12'h000;
      20'h01e6d: out <= 12'h000;
      20'h01e6e: out <= 12'h000;
      20'h01e6f: out <= 12'h000;
      20'h01e70: out <= 12'h000;
      20'h01e71: out <= 12'h000;
      20'h01e72: out <= 12'h000;
      20'h01e73: out <= 12'h000;
      20'h01e74: out <= 12'h000;
      20'h01e75: out <= 12'h000;
      20'h01e76: out <= 12'h000;
      20'h01e77: out <= 12'h000;
      20'h01e78: out <= 12'h000;
      20'h01e79: out <= 12'h000;
      20'h01e7a: out <= 12'h000;
      20'h01e7b: out <= 12'h000;
      20'h01e7c: out <= 12'h000;
      20'h01e7d: out <= 12'h000;
      20'h01e7e: out <= 12'h000;
      20'h01e7f: out <= 12'h000;
      20'h01e80: out <= 12'h000;
      20'h01e81: out <= 12'h000;
      20'h01e82: out <= 12'h000;
      20'h01e83: out <= 12'h000;
      20'h01e84: out <= 12'h000;
      20'h01e85: out <= 12'h000;
      20'h01e86: out <= 12'h000;
      20'h01e87: out <= 12'h000;
      20'h01e88: out <= 12'h000;
      20'h01e89: out <= 12'h000;
      20'h01e8a: out <= 12'h000;
      20'h01e8b: out <= 12'h000;
      20'h01e8c: out <= 12'h000;
      20'h01e8d: out <= 12'h000;
      20'h01e8e: out <= 12'h000;
      20'h01e8f: out <= 12'h000;
      20'h01e90: out <= 12'h000;
      20'h01e91: out <= 12'h000;
      20'h01e92: out <= 12'h000;
      20'h01e93: out <= 12'h000;
      20'h01e94: out <= 12'h000;
      20'h01e95: out <= 12'h000;
      20'h01e96: out <= 12'h000;
      20'h01e97: out <= 12'h000;
      20'h01e98: out <= 12'h000;
      20'h01e99: out <= 12'h000;
      20'h01e9a: out <= 12'h000;
      20'h01e9b: out <= 12'h000;
      20'h01e9c: out <= 12'h000;
      20'h01e9d: out <= 12'h000;
      20'h01e9e: out <= 12'h000;
      20'h01e9f: out <= 12'h000;
      20'h01ea0: out <= 12'h000;
      20'h01ea1: out <= 12'h6af;
      20'h01ea2: out <= 12'hfff;
      20'h01ea3: out <= 12'h6af;
      20'h01ea4: out <= 12'h16d;
      20'h01ea5: out <= 12'h16d;
      20'h01ea6: out <= 12'h16d;
      20'h01ea7: out <= 12'h16d;
      20'h01ea8: out <= 12'h16d;
      20'h01ea9: out <= 12'h6af;
      20'h01eaa: out <= 12'hfff;
      20'h01eab: out <= 12'hfff;
      20'h01eac: out <= 12'h6af;
      20'h01ead: out <= 12'h000;
      20'h01eae: out <= 12'h000;
      20'h01eaf: out <= 12'h000;
      20'h01eb0: out <= 12'h222;
      20'h01eb1: out <= 12'h6af;
      20'h01eb2: out <= 12'hfff;
      20'h01eb3: out <= 12'h6af;
      20'h01eb4: out <= 12'hfff;
      20'h01eb5: out <= 12'hfff;
      20'h01eb6: out <= 12'hfff;
      20'h01eb7: out <= 12'hfff;
      20'h01eb8: out <= 12'hfff;
      20'h01eb9: out <= 12'h6af;
      20'h01eba: out <= 12'h16d;
      20'h01ebb: out <= 12'hfff;
      20'h01ebc: out <= 12'h6af;
      20'h01ebd: out <= 12'h222;
      20'h01ebe: out <= 12'h222;
      20'h01ebf: out <= 12'h222;
      20'h01ec0: out <= 12'h000;
      20'h01ec1: out <= 12'h6af;
      20'h01ec2: out <= 12'hfff;
      20'h01ec3: out <= 12'h6af;
      20'h01ec4: out <= 12'h16d;
      20'h01ec5: out <= 12'h16d;
      20'h01ec6: out <= 12'h6af;
      20'h01ec7: out <= 12'hfff;
      20'h01ec8: out <= 12'hfff;
      20'h01ec9: out <= 12'hfff;
      20'h01eca: out <= 12'h6af;
      20'h01ecb: out <= 12'h16d;
      20'h01ecc: out <= 12'h16d;
      20'h01ecd: out <= 12'h6af;
      20'h01ece: out <= 12'hfff;
      20'h01ecf: out <= 12'h6af;
      20'h01ed0: out <= 12'h222;
      20'h01ed1: out <= 12'h6af;
      20'h01ed2: out <= 12'h16d;
      20'h01ed3: out <= 12'h6af;
      20'h01ed4: out <= 12'hfff;
      20'h01ed5: out <= 12'hfff;
      20'h01ed6: out <= 12'h6af;
      20'h01ed7: out <= 12'hfff;
      20'h01ed8: out <= 12'hfff;
      20'h01ed9: out <= 12'hfff;
      20'h01eda: out <= 12'h6af;
      20'h01edb: out <= 12'hfff;
      20'h01edc: out <= 12'hfff;
      20'h01edd: out <= 12'h6af;
      20'h01ede: out <= 12'h16d;
      20'h01edf: out <= 12'h6af;
      20'h01ee0: out <= 12'h000;
      20'h01ee1: out <= 12'h000;
      20'h01ee2: out <= 12'h000;
      20'h01ee3: out <= 12'h6af;
      20'h01ee4: out <= 12'hfff;
      20'h01ee5: out <= 12'hfff;
      20'h01ee6: out <= 12'h6af;
      20'h01ee7: out <= 12'h16d;
      20'h01ee8: out <= 12'h16d;
      20'h01ee9: out <= 12'h16d;
      20'h01eea: out <= 12'h16d;
      20'h01eeb: out <= 12'h16d;
      20'h01eec: out <= 12'h6af;
      20'h01eed: out <= 12'hfff;
      20'h01eee: out <= 12'h6af;
      20'h01eef: out <= 12'h000;
      20'h01ef0: out <= 12'h222;
      20'h01ef1: out <= 12'h222;
      20'h01ef2: out <= 12'h222;
      20'h01ef3: out <= 12'h6af;
      20'h01ef4: out <= 12'hfff;
      20'h01ef5: out <= 12'h16d;
      20'h01ef6: out <= 12'h6af;
      20'h01ef7: out <= 12'hfff;
      20'h01ef8: out <= 12'hfff;
      20'h01ef9: out <= 12'hfff;
      20'h01efa: out <= 12'hfff;
      20'h01efb: out <= 12'hfff;
      20'h01efc: out <= 12'h6af;
      20'h01efd: out <= 12'hfff;
      20'h01efe: out <= 12'h6af;
      20'h01eff: out <= 12'h222;
      20'h01f00: out <= 12'h000;
      20'h01f01: out <= 12'h6af;
      20'h01f02: out <= 12'h16d;
      20'h01f03: out <= 12'h6af;
      20'h01f04: out <= 12'h000;
      20'h01f05: out <= 12'h000;
      20'h01f06: out <= 12'hfff;
      20'h01f07: out <= 12'hfff;
      20'h01f08: out <= 12'hfff;
      20'h01f09: out <= 12'hfff;
      20'h01f0a: out <= 12'hfff;
      20'h01f0b: out <= 12'h000;
      20'h01f0c: out <= 12'h000;
      20'h01f0d: out <= 12'h6af;
      20'h01f0e: out <= 12'h16d;
      20'h01f0f: out <= 12'h6af;
      20'h01f10: out <= 12'h222;
      20'h01f11: out <= 12'h6af;
      20'h01f12: out <= 12'h16d;
      20'h01f13: out <= 12'h6af;
      20'h01f14: out <= 12'h222;
      20'h01f15: out <= 12'h222;
      20'h01f16: out <= 12'h16d;
      20'h01f17: out <= 12'h16d;
      20'h01f18: out <= 12'h16d;
      20'h01f19: out <= 12'h16d;
      20'h01f1a: out <= 12'h16d;
      20'h01f1b: out <= 12'h222;
      20'h01f1c: out <= 12'h222;
      20'h01f1d: out <= 12'h6af;
      20'h01f1e: out <= 12'h16d;
      20'h01f1f: out <= 12'h6af;
      20'h01f20: out <= 12'h603;
      20'h01f21: out <= 12'h603;
      20'h01f22: out <= 12'h603;
      20'h01f23: out <= 12'h603;
      20'h01f24: out <= 12'hfff;
      20'h01f25: out <= 12'hbbb;
      20'h01f26: out <= 12'h666;
      20'h01f27: out <= 12'hfff;
      20'h01f28: out <= 12'hfff;
      20'h01f29: out <= 12'hbbb;
      20'h01f2a: out <= 12'h666;
      20'h01f2b: out <= 12'h666;
      20'h01f2c: out <= 12'hfff;
      20'h01f2d: out <= 12'hbbb;
      20'h01f2e: out <= 12'h666;
      20'h01f2f: out <= 12'hfff;
      20'h01f30: out <= 12'hfff;
      20'h01f31: out <= 12'hbbb;
      20'h01f32: out <= 12'h666;
      20'h01f33: out <= 12'h666;
      20'h01f34: out <= 12'h000;
      20'h01f35: out <= 12'h000;
      20'h01f36: out <= 12'h000;
      20'h01f37: out <= 12'h000;
      20'h01f38: out <= 12'h000;
      20'h01f39: out <= 12'h000;
      20'h01f3a: out <= 12'h000;
      20'h01f3b: out <= 12'h000;
      20'h01f3c: out <= 12'hfff;
      20'h01f3d: out <= 12'hbbb;
      20'h01f3e: out <= 12'h666;
      20'h01f3f: out <= 12'hfff;
      20'h01f40: out <= 12'hfff;
      20'h01f41: out <= 12'hbbb;
      20'h01f42: out <= 12'h666;
      20'h01f43: out <= 12'h666;
      20'h01f44: out <= 12'hfff;
      20'h01f45: out <= 12'hbbb;
      20'h01f46: out <= 12'h666;
      20'h01f47: out <= 12'hfff;
      20'h01f48: out <= 12'hfff;
      20'h01f49: out <= 12'hbbb;
      20'h01f4a: out <= 12'h666;
      20'h01f4b: out <= 12'h666;
      20'h01f4c: out <= 12'hfff;
      20'h01f4d: out <= 12'hbbb;
      20'h01f4e: out <= 12'h666;
      20'h01f4f: out <= 12'hfff;
      20'h01f50: out <= 12'hfff;
      20'h01f51: out <= 12'hbbb;
      20'h01f52: out <= 12'h666;
      20'h01f53: out <= 12'h666;
      20'h01f54: out <= 12'hfff;
      20'h01f55: out <= 12'hbbb;
      20'h01f56: out <= 12'h666;
      20'h01f57: out <= 12'hfff;
      20'h01f58: out <= 12'hfff;
      20'h01f59: out <= 12'hbbb;
      20'h01f5a: out <= 12'h666;
      20'h01f5b: out <= 12'h666;
      20'h01f5c: out <= 12'h000;
      20'h01f5d: out <= 12'h000;
      20'h01f5e: out <= 12'h000;
      20'h01f5f: out <= 12'h000;
      20'h01f60: out <= 12'h000;
      20'h01f61: out <= 12'h000;
      20'h01f62: out <= 12'h000;
      20'h01f63: out <= 12'h000;
      20'h01f64: out <= 12'h000;
      20'h01f65: out <= 12'h000;
      20'h01f66: out <= 12'h000;
      20'h01f67: out <= 12'h000;
      20'h01f68: out <= 12'h000;
      20'h01f69: out <= 12'h000;
      20'h01f6a: out <= 12'h000;
      20'h01f6b: out <= 12'h000;
      20'h01f6c: out <= 12'h000;
      20'h01f6d: out <= 12'h000;
      20'h01f6e: out <= 12'h000;
      20'h01f6f: out <= 12'h000;
      20'h01f70: out <= 12'h000;
      20'h01f71: out <= 12'h000;
      20'h01f72: out <= 12'h000;
      20'h01f73: out <= 12'h000;
      20'h01f74: out <= 12'h603;
      20'h01f75: out <= 12'h603;
      20'h01f76: out <= 12'h603;
      20'h01f77: out <= 12'h603;
      20'h01f78: out <= 12'hee9;
      20'h01f79: out <= 12'hf87;
      20'h01f7a: out <= 12'hee9;
      20'h01f7b: out <= 12'hf87;
      20'h01f7c: out <= 12'hf87;
      20'h01f7d: out <= 12'hb27;
      20'h01f7e: out <= 12'hf87;
      20'h01f7f: out <= 12'hb27;
      20'h01f80: out <= 12'h000;
      20'h01f81: out <= 12'h000;
      20'h01f82: out <= 12'h000;
      20'h01f83: out <= 12'h000;
      20'h01f84: out <= 12'h000;
      20'h01f85: out <= 12'h000;
      20'h01f86: out <= 12'h000;
      20'h01f87: out <= 12'h000;
      20'h01f88: out <= 12'h000;
      20'h01f89: out <= 12'h000;
      20'h01f8a: out <= 12'h000;
      20'h01f8b: out <= 12'h000;
      20'h01f8c: out <= 12'h000;
      20'h01f8d: out <= 12'h000;
      20'h01f8e: out <= 12'h000;
      20'h01f8f: out <= 12'h000;
      20'h01f90: out <= 12'h000;
      20'h01f91: out <= 12'h000;
      20'h01f92: out <= 12'h000;
      20'h01f93: out <= 12'h000;
      20'h01f94: out <= 12'h000;
      20'h01f95: out <= 12'h000;
      20'h01f96: out <= 12'h000;
      20'h01f97: out <= 12'h000;
      20'h01f98: out <= 12'h000;
      20'h01f99: out <= 12'h000;
      20'h01f9a: out <= 12'h000;
      20'h01f9b: out <= 12'h000;
      20'h01f9c: out <= 12'h000;
      20'h01f9d: out <= 12'h000;
      20'h01f9e: out <= 12'h000;
      20'h01f9f: out <= 12'h000;
      20'h01fa0: out <= 12'h000;
      20'h01fa1: out <= 12'h000;
      20'h01fa2: out <= 12'h000;
      20'h01fa3: out <= 12'h000;
      20'h01fa4: out <= 12'h000;
      20'h01fa5: out <= 12'h000;
      20'h01fa6: out <= 12'h000;
      20'h01fa7: out <= 12'h000;
      20'h01fa8: out <= 12'h000;
      20'h01fa9: out <= 12'h000;
      20'h01faa: out <= 12'h000;
      20'h01fab: out <= 12'h000;
      20'h01fac: out <= 12'h000;
      20'h01fad: out <= 12'h000;
      20'h01fae: out <= 12'h000;
      20'h01faf: out <= 12'h000;
      20'h01fb0: out <= 12'h000;
      20'h01fb1: out <= 12'h000;
      20'h01fb2: out <= 12'h000;
      20'h01fb3: out <= 12'h000;
      20'h01fb4: out <= 12'h000;
      20'h01fb5: out <= 12'h000;
      20'h01fb6: out <= 12'h000;
      20'h01fb7: out <= 12'h000;
      20'h01fb8: out <= 12'h000;
      20'h01fb9: out <= 12'h16d;
      20'h01fba: out <= 12'hfff;
      20'h01fbb: out <= 12'hfff;
      20'h01fbc: out <= 12'h6af;
      20'h01fbd: out <= 12'h6af;
      20'h01fbe: out <= 12'h6af;
      20'h01fbf: out <= 12'h6af;
      20'h01fc0: out <= 12'h6af;
      20'h01fc1: out <= 12'hfff;
      20'h01fc2: out <= 12'h16d;
      20'h01fc3: out <= 12'hfff;
      20'h01fc4: out <= 12'h16d;
      20'h01fc5: out <= 12'h000;
      20'h01fc6: out <= 12'h000;
      20'h01fc7: out <= 12'h000;
      20'h01fc8: out <= 12'h222;
      20'h01fc9: out <= 12'h16d;
      20'h01fca: out <= 12'hfff;
      20'h01fcb: out <= 12'h16d;
      20'h01fcc: out <= 12'h6af;
      20'h01fcd: out <= 12'h6af;
      20'h01fce: out <= 12'h6af;
      20'h01fcf: out <= 12'h6af;
      20'h01fd0: out <= 12'h6af;
      20'h01fd1: out <= 12'h16d;
      20'h01fd2: out <= 12'h16d;
      20'h01fd3: out <= 12'hfff;
      20'h01fd4: out <= 12'h16d;
      20'h01fd5: out <= 12'h222;
      20'h01fd6: out <= 12'h222;
      20'h01fd7: out <= 12'h222;
      20'h01fd8: out <= 12'h000;
      20'h01fd9: out <= 12'hfff;
      20'h01fda: out <= 12'hfff;
      20'h01fdb: out <= 12'hfff;
      20'h01fdc: out <= 12'h6af;
      20'h01fdd: out <= 12'h6af;
      20'h01fde: out <= 12'h16d;
      20'h01fdf: out <= 12'h16d;
      20'h01fe0: out <= 12'h16d;
      20'h01fe1: out <= 12'h16d;
      20'h01fe2: out <= 12'h16d;
      20'h01fe3: out <= 12'h6af;
      20'h01fe4: out <= 12'h6af;
      20'h01fe5: out <= 12'hfff;
      20'h01fe6: out <= 12'hfff;
      20'h01fe7: out <= 12'hfff;
      20'h01fe8: out <= 12'h222;
      20'h01fe9: out <= 12'hfff;
      20'h01fea: out <= 12'hfff;
      20'h01feb: out <= 12'hfff;
      20'h01fec: out <= 12'h6af;
      20'h01fed: out <= 12'h6af;
      20'h01fee: out <= 12'hfff;
      20'h01fef: out <= 12'hfff;
      20'h01ff0: out <= 12'hfff;
      20'h01ff1: out <= 12'hfff;
      20'h01ff2: out <= 12'hfff;
      20'h01ff3: out <= 12'h6af;
      20'h01ff4: out <= 12'h6af;
      20'h01ff5: out <= 12'hfff;
      20'h01ff6: out <= 12'hfff;
      20'h01ff7: out <= 12'hfff;
      20'h01ff8: out <= 12'h000;
      20'h01ff9: out <= 12'h000;
      20'h01ffa: out <= 12'h000;
      20'h01ffb: out <= 12'h16d;
      20'h01ffc: out <= 12'hfff;
      20'h01ffd: out <= 12'h16d;
      20'h01ffe: out <= 12'hfff;
      20'h01fff: out <= 12'h6af;
      20'h02000: out <= 12'h6af;
      20'h02001: out <= 12'h6af;
      20'h02002: out <= 12'h6af;
      20'h02003: out <= 12'h6af;
      20'h02004: out <= 12'hfff;
      20'h02005: out <= 12'hfff;
      20'h02006: out <= 12'h16d;
      20'h02007: out <= 12'h000;
      20'h02008: out <= 12'h222;
      20'h02009: out <= 12'h222;
      20'h0200a: out <= 12'h222;
      20'h0200b: out <= 12'h16d;
      20'h0200c: out <= 12'hfff;
      20'h0200d: out <= 12'h16d;
      20'h0200e: out <= 12'h16d;
      20'h0200f: out <= 12'h6af;
      20'h02010: out <= 12'h6af;
      20'h02011: out <= 12'h6af;
      20'h02012: out <= 12'h6af;
      20'h02013: out <= 12'h6af;
      20'h02014: out <= 12'h16d;
      20'h02015: out <= 12'hfff;
      20'h02016: out <= 12'h16d;
      20'h02017: out <= 12'h222;
      20'h02018: out <= 12'h000;
      20'h02019: out <= 12'h000;
      20'h0201a: out <= 12'h000;
      20'h0201b: out <= 12'h000;
      20'h0201c: out <= 12'h000;
      20'h0201d: out <= 12'h000;
      20'h0201e: out <= 12'h000;
      20'h0201f: out <= 12'h16d;
      20'h02020: out <= 12'hfff;
      20'h02021: out <= 12'h16d;
      20'h02022: out <= 12'h000;
      20'h02023: out <= 12'h000;
      20'h02024: out <= 12'h000;
      20'h02025: out <= 12'h000;
      20'h02026: out <= 12'h000;
      20'h02027: out <= 12'h000;
      20'h02028: out <= 12'h222;
      20'h02029: out <= 12'h222;
      20'h0202a: out <= 12'h222;
      20'h0202b: out <= 12'h222;
      20'h0202c: out <= 12'h222;
      20'h0202d: out <= 12'h222;
      20'h0202e: out <= 12'h222;
      20'h0202f: out <= 12'h16d;
      20'h02030: out <= 12'hfff;
      20'h02031: out <= 12'h16d;
      20'h02032: out <= 12'h222;
      20'h02033: out <= 12'h222;
      20'h02034: out <= 12'h222;
      20'h02035: out <= 12'h222;
      20'h02036: out <= 12'h222;
      20'h02037: out <= 12'h222;
      20'h02038: out <= 12'h603;
      20'h02039: out <= 12'h603;
      20'h0203a: out <= 12'h603;
      20'h0203b: out <= 12'h603;
      20'h0203c: out <= 12'hfff;
      20'h0203d: out <= 12'hbbb;
      20'h0203e: out <= 12'hbbb;
      20'h0203f: out <= 12'hbbb;
      20'h02040: out <= 12'hbbb;
      20'h02041: out <= 12'hbbb;
      20'h02042: out <= 12'h666;
      20'h02043: out <= 12'h666;
      20'h02044: out <= 12'hfff;
      20'h02045: out <= 12'hbbb;
      20'h02046: out <= 12'hbbb;
      20'h02047: out <= 12'hbbb;
      20'h02048: out <= 12'hbbb;
      20'h02049: out <= 12'hbbb;
      20'h0204a: out <= 12'h666;
      20'h0204b: out <= 12'h666;
      20'h0204c: out <= 12'h000;
      20'h0204d: out <= 12'h000;
      20'h0204e: out <= 12'h000;
      20'h0204f: out <= 12'h000;
      20'h02050: out <= 12'h000;
      20'h02051: out <= 12'h000;
      20'h02052: out <= 12'h000;
      20'h02053: out <= 12'h000;
      20'h02054: out <= 12'hfff;
      20'h02055: out <= 12'hbbb;
      20'h02056: out <= 12'hbbb;
      20'h02057: out <= 12'hbbb;
      20'h02058: out <= 12'hbbb;
      20'h02059: out <= 12'hbbb;
      20'h0205a: out <= 12'h666;
      20'h0205b: out <= 12'h666;
      20'h0205c: out <= 12'hfff;
      20'h0205d: out <= 12'hbbb;
      20'h0205e: out <= 12'hbbb;
      20'h0205f: out <= 12'hbbb;
      20'h02060: out <= 12'hbbb;
      20'h02061: out <= 12'hbbb;
      20'h02062: out <= 12'h666;
      20'h02063: out <= 12'h666;
      20'h02064: out <= 12'hfff;
      20'h02065: out <= 12'hbbb;
      20'h02066: out <= 12'hbbb;
      20'h02067: out <= 12'hbbb;
      20'h02068: out <= 12'hbbb;
      20'h02069: out <= 12'hbbb;
      20'h0206a: out <= 12'h666;
      20'h0206b: out <= 12'h666;
      20'h0206c: out <= 12'hfff;
      20'h0206d: out <= 12'hbbb;
      20'h0206e: out <= 12'hbbb;
      20'h0206f: out <= 12'hbbb;
      20'h02070: out <= 12'hbbb;
      20'h02071: out <= 12'hbbb;
      20'h02072: out <= 12'h666;
      20'h02073: out <= 12'h666;
      20'h02074: out <= 12'h000;
      20'h02075: out <= 12'h000;
      20'h02076: out <= 12'h000;
      20'h02077: out <= 12'h000;
      20'h02078: out <= 12'h000;
      20'h02079: out <= 12'h000;
      20'h0207a: out <= 12'h000;
      20'h0207b: out <= 12'h000;
      20'h0207c: out <= 12'h000;
      20'h0207d: out <= 12'h000;
      20'h0207e: out <= 12'h000;
      20'h0207f: out <= 12'h000;
      20'h02080: out <= 12'h000;
      20'h02081: out <= 12'h000;
      20'h02082: out <= 12'h000;
      20'h02083: out <= 12'h000;
      20'h02084: out <= 12'h000;
      20'h02085: out <= 12'h000;
      20'h02086: out <= 12'h000;
      20'h02087: out <= 12'h000;
      20'h02088: out <= 12'h000;
      20'h02089: out <= 12'h000;
      20'h0208a: out <= 12'h000;
      20'h0208b: out <= 12'h000;
      20'h0208c: out <= 12'h603;
      20'h0208d: out <= 12'h603;
      20'h0208e: out <= 12'h603;
      20'h0208f: out <= 12'h603;
      20'h02090: out <= 12'hee9;
      20'h02091: out <= 12'hf87;
      20'h02092: out <= 12'hee9;
      20'h02093: out <= 12'hb27;
      20'h02094: out <= 12'hb27;
      20'h02095: out <= 12'hb27;
      20'h02096: out <= 12'hf87;
      20'h02097: out <= 12'hb27;
      20'h02098: out <= 12'h000;
      20'h02099: out <= 12'h000;
      20'h0209a: out <= 12'h000;
      20'h0209b: out <= 12'h000;
      20'h0209c: out <= 12'h000;
      20'h0209d: out <= 12'h000;
      20'h0209e: out <= 12'h000;
      20'h0209f: out <= 12'h000;
      20'h020a0: out <= 12'h000;
      20'h020a1: out <= 12'h000;
      20'h020a2: out <= 12'h000;
      20'h020a3: out <= 12'h000;
      20'h020a4: out <= 12'h000;
      20'h020a5: out <= 12'h000;
      20'h020a6: out <= 12'h000;
      20'h020a7: out <= 12'h000;
      20'h020a8: out <= 12'h000;
      20'h020a9: out <= 12'h000;
      20'h020aa: out <= 12'h000;
      20'h020ab: out <= 12'h000;
      20'h020ac: out <= 12'h000;
      20'h020ad: out <= 12'h000;
      20'h020ae: out <= 12'h000;
      20'h020af: out <= 12'h000;
      20'h020b0: out <= 12'h000;
      20'h020b1: out <= 12'h000;
      20'h020b2: out <= 12'h000;
      20'h020b3: out <= 12'h000;
      20'h020b4: out <= 12'h000;
      20'h020b5: out <= 12'h000;
      20'h020b6: out <= 12'h000;
      20'h020b7: out <= 12'h000;
      20'h020b8: out <= 12'h000;
      20'h020b9: out <= 12'h000;
      20'h020ba: out <= 12'h000;
      20'h020bb: out <= 12'h000;
      20'h020bc: out <= 12'h000;
      20'h020bd: out <= 12'h000;
      20'h020be: out <= 12'h000;
      20'h020bf: out <= 12'h000;
      20'h020c0: out <= 12'h000;
      20'h020c1: out <= 12'h000;
      20'h020c2: out <= 12'h000;
      20'h020c3: out <= 12'h000;
      20'h020c4: out <= 12'h000;
      20'h020c5: out <= 12'h000;
      20'h020c6: out <= 12'h000;
      20'h020c7: out <= 12'h000;
      20'h020c8: out <= 12'h000;
      20'h020c9: out <= 12'h000;
      20'h020ca: out <= 12'h000;
      20'h020cb: out <= 12'h000;
      20'h020cc: out <= 12'h000;
      20'h020cd: out <= 12'h000;
      20'h020ce: out <= 12'h000;
      20'h020cf: out <= 12'h000;
      20'h020d0: out <= 12'h000;
      20'h020d1: out <= 12'h6af;
      20'h020d2: out <= 12'hfff;
      20'h020d3: out <= 12'h6af;
      20'h020d4: out <= 12'hfff;
      20'h020d5: out <= 12'hfff;
      20'h020d6: out <= 12'hfff;
      20'h020d7: out <= 12'hfff;
      20'h020d8: out <= 12'hfff;
      20'h020d9: out <= 12'h6af;
      20'h020da: out <= 12'h6af;
      20'h020db: out <= 12'hfff;
      20'h020dc: out <= 12'h6af;
      20'h020dd: out <= 12'h000;
      20'h020de: out <= 12'h000;
      20'h020df: out <= 12'h000;
      20'h020e0: out <= 12'h222;
      20'h020e1: out <= 12'h6af;
      20'h020e2: out <= 12'hfff;
      20'h020e3: out <= 12'h6af;
      20'h020e4: out <= 12'h16d;
      20'h020e5: out <= 12'h16d;
      20'h020e6: out <= 12'h16d;
      20'h020e7: out <= 12'h16d;
      20'h020e8: out <= 12'h16d;
      20'h020e9: out <= 12'h6af;
      20'h020ea: out <= 12'h6af;
      20'h020eb: out <= 12'hfff;
      20'h020ec: out <= 12'h6af;
      20'h020ed: out <= 12'h222;
      20'h020ee: out <= 12'h222;
      20'h020ef: out <= 12'h222;
      20'h020f0: out <= 12'h000;
      20'h020f1: out <= 12'h6af;
      20'h020f2: out <= 12'h16d;
      20'h020f3: out <= 12'h6af;
      20'h020f4: out <= 12'hfff;
      20'h020f5: out <= 12'hfff;
      20'h020f6: out <= 12'h6af;
      20'h020f7: out <= 12'h6af;
      20'h020f8: out <= 12'h6af;
      20'h020f9: out <= 12'h6af;
      20'h020fa: out <= 12'h6af;
      20'h020fb: out <= 12'hfff;
      20'h020fc: out <= 12'hfff;
      20'h020fd: out <= 12'h6af;
      20'h020fe: out <= 12'h16d;
      20'h020ff: out <= 12'h6af;
      20'h02100: out <= 12'h222;
      20'h02101: out <= 12'h6af;
      20'h02102: out <= 12'h16d;
      20'h02103: out <= 12'h6af;
      20'h02104: out <= 12'h16d;
      20'h02105: out <= 12'h16d;
      20'h02106: out <= 12'h6af;
      20'h02107: out <= 12'h6af;
      20'h02108: out <= 12'h6af;
      20'h02109: out <= 12'h6af;
      20'h0210a: out <= 12'h6af;
      20'h0210b: out <= 12'h16d;
      20'h0210c: out <= 12'h16d;
      20'h0210d: out <= 12'h6af;
      20'h0210e: out <= 12'h16d;
      20'h0210f: out <= 12'h6af;
      20'h02110: out <= 12'h000;
      20'h02111: out <= 12'h000;
      20'h02112: out <= 12'h000;
      20'h02113: out <= 12'h6af;
      20'h02114: out <= 12'hfff;
      20'h02115: out <= 12'h6af;
      20'h02116: out <= 12'h6af;
      20'h02117: out <= 12'hfff;
      20'h02118: out <= 12'hfff;
      20'h02119: out <= 12'hfff;
      20'h0211a: out <= 12'hfff;
      20'h0211b: out <= 12'hfff;
      20'h0211c: out <= 12'h6af;
      20'h0211d: out <= 12'hfff;
      20'h0211e: out <= 12'h6af;
      20'h0211f: out <= 12'h000;
      20'h02120: out <= 12'h222;
      20'h02121: out <= 12'h222;
      20'h02122: out <= 12'h222;
      20'h02123: out <= 12'h6af;
      20'h02124: out <= 12'hfff;
      20'h02125: out <= 12'h6af;
      20'h02126: out <= 12'h6af;
      20'h02127: out <= 12'h16d;
      20'h02128: out <= 12'h16d;
      20'h02129: out <= 12'h16d;
      20'h0212a: out <= 12'h16d;
      20'h0212b: out <= 12'h16d;
      20'h0212c: out <= 12'h6af;
      20'h0212d: out <= 12'hfff;
      20'h0212e: out <= 12'h6af;
      20'h0212f: out <= 12'h222;
      20'h02130: out <= 12'h000;
      20'h02131: out <= 12'h000;
      20'h02132: out <= 12'h000;
      20'h02133: out <= 12'h000;
      20'h02134: out <= 12'h000;
      20'h02135: out <= 12'h000;
      20'h02136: out <= 12'h000;
      20'h02137: out <= 12'h16d;
      20'h02138: out <= 12'hfff;
      20'h02139: out <= 12'h16d;
      20'h0213a: out <= 12'h000;
      20'h0213b: out <= 12'h000;
      20'h0213c: out <= 12'h000;
      20'h0213d: out <= 12'h000;
      20'h0213e: out <= 12'h000;
      20'h0213f: out <= 12'h000;
      20'h02140: out <= 12'h222;
      20'h02141: out <= 12'h222;
      20'h02142: out <= 12'h222;
      20'h02143: out <= 12'h222;
      20'h02144: out <= 12'h222;
      20'h02145: out <= 12'h222;
      20'h02146: out <= 12'h222;
      20'h02147: out <= 12'h16d;
      20'h02148: out <= 12'hfff;
      20'h02149: out <= 12'h16d;
      20'h0214a: out <= 12'h222;
      20'h0214b: out <= 12'h222;
      20'h0214c: out <= 12'h222;
      20'h0214d: out <= 12'h222;
      20'h0214e: out <= 12'h222;
      20'h0214f: out <= 12'h222;
      20'h02150: out <= 12'h603;
      20'h02151: out <= 12'h603;
      20'h02152: out <= 12'h603;
      20'h02153: out <= 12'h603;
      20'h02154: out <= 12'hfff;
      20'h02155: out <= 12'h666;
      20'h02156: out <= 12'h666;
      20'h02157: out <= 12'h666;
      20'h02158: out <= 12'h666;
      20'h02159: out <= 12'h666;
      20'h0215a: out <= 12'h666;
      20'h0215b: out <= 12'h666;
      20'h0215c: out <= 12'hfff;
      20'h0215d: out <= 12'h666;
      20'h0215e: out <= 12'h666;
      20'h0215f: out <= 12'h666;
      20'h02160: out <= 12'h666;
      20'h02161: out <= 12'h666;
      20'h02162: out <= 12'h666;
      20'h02163: out <= 12'h666;
      20'h02164: out <= 12'h000;
      20'h02165: out <= 12'h000;
      20'h02166: out <= 12'h000;
      20'h02167: out <= 12'h000;
      20'h02168: out <= 12'h000;
      20'h02169: out <= 12'h000;
      20'h0216a: out <= 12'h000;
      20'h0216b: out <= 12'h000;
      20'h0216c: out <= 12'hfff;
      20'h0216d: out <= 12'h666;
      20'h0216e: out <= 12'h666;
      20'h0216f: out <= 12'h666;
      20'h02170: out <= 12'h666;
      20'h02171: out <= 12'h666;
      20'h02172: out <= 12'h666;
      20'h02173: out <= 12'h666;
      20'h02174: out <= 12'hfff;
      20'h02175: out <= 12'h666;
      20'h02176: out <= 12'h666;
      20'h02177: out <= 12'h666;
      20'h02178: out <= 12'h666;
      20'h02179: out <= 12'h666;
      20'h0217a: out <= 12'h666;
      20'h0217b: out <= 12'h666;
      20'h0217c: out <= 12'hfff;
      20'h0217d: out <= 12'h666;
      20'h0217e: out <= 12'h666;
      20'h0217f: out <= 12'h666;
      20'h02180: out <= 12'h666;
      20'h02181: out <= 12'h666;
      20'h02182: out <= 12'h666;
      20'h02183: out <= 12'h666;
      20'h02184: out <= 12'hfff;
      20'h02185: out <= 12'h666;
      20'h02186: out <= 12'h666;
      20'h02187: out <= 12'h666;
      20'h02188: out <= 12'h666;
      20'h02189: out <= 12'h666;
      20'h0218a: out <= 12'h666;
      20'h0218b: out <= 12'h666;
      20'h0218c: out <= 12'h000;
      20'h0218d: out <= 12'h000;
      20'h0218e: out <= 12'h000;
      20'h0218f: out <= 12'h000;
      20'h02190: out <= 12'h000;
      20'h02191: out <= 12'h000;
      20'h02192: out <= 12'h000;
      20'h02193: out <= 12'h000;
      20'h02194: out <= 12'h000;
      20'h02195: out <= 12'h000;
      20'h02196: out <= 12'h000;
      20'h02197: out <= 12'h000;
      20'h02198: out <= 12'h000;
      20'h02199: out <= 12'h000;
      20'h0219a: out <= 12'h000;
      20'h0219b: out <= 12'h000;
      20'h0219c: out <= 12'h000;
      20'h0219d: out <= 12'h000;
      20'h0219e: out <= 12'h000;
      20'h0219f: out <= 12'h000;
      20'h021a0: out <= 12'h000;
      20'h021a1: out <= 12'h000;
      20'h021a2: out <= 12'h000;
      20'h021a3: out <= 12'h000;
      20'h021a4: out <= 12'h603;
      20'h021a5: out <= 12'h603;
      20'h021a6: out <= 12'h603;
      20'h021a7: out <= 12'h603;
      20'h021a8: out <= 12'hee9;
      20'h021a9: out <= 12'hf87;
      20'h021aa: out <= 12'hf87;
      20'h021ab: out <= 12'hf87;
      20'h021ac: out <= 12'hf87;
      20'h021ad: out <= 12'hf87;
      20'h021ae: out <= 12'hf87;
      20'h021af: out <= 12'hb27;
      20'h021b0: out <= 12'h000;
      20'h021b1: out <= 12'h000;
      20'h021b2: out <= 12'h000;
      20'h021b3: out <= 12'h000;
      20'h021b4: out <= 12'h000;
      20'h021b5: out <= 12'h000;
      20'h021b6: out <= 12'h000;
      20'h021b7: out <= 12'h000;
      20'h021b8: out <= 12'h000;
      20'h021b9: out <= 12'h000;
      20'h021ba: out <= 12'h000;
      20'h021bb: out <= 12'h000;
      20'h021bc: out <= 12'h000;
      20'h021bd: out <= 12'h000;
      20'h021be: out <= 12'h000;
      20'h021bf: out <= 12'h000;
      20'h021c0: out <= 12'h000;
      20'h021c1: out <= 12'h000;
      20'h021c2: out <= 12'h000;
      20'h021c3: out <= 12'h000;
      20'h021c4: out <= 12'h000;
      20'h021c5: out <= 12'h000;
      20'h021c6: out <= 12'h000;
      20'h021c7: out <= 12'h000;
      20'h021c8: out <= 12'h000;
      20'h021c9: out <= 12'h000;
      20'h021ca: out <= 12'h000;
      20'h021cb: out <= 12'h000;
      20'h021cc: out <= 12'h000;
      20'h021cd: out <= 12'h000;
      20'h021ce: out <= 12'h000;
      20'h021cf: out <= 12'h000;
      20'h021d0: out <= 12'h000;
      20'h021d1: out <= 12'h000;
      20'h021d2: out <= 12'h000;
      20'h021d3: out <= 12'h000;
      20'h021d4: out <= 12'h000;
      20'h021d5: out <= 12'h000;
      20'h021d6: out <= 12'h000;
      20'h021d7: out <= 12'h000;
      20'h021d8: out <= 12'h000;
      20'h021d9: out <= 12'h000;
      20'h021da: out <= 12'h000;
      20'h021db: out <= 12'h000;
      20'h021dc: out <= 12'h000;
      20'h021dd: out <= 12'h000;
      20'h021de: out <= 12'h000;
      20'h021df: out <= 12'h000;
      20'h021e0: out <= 12'h000;
      20'h021e1: out <= 12'h000;
      20'h021e2: out <= 12'h000;
      20'h021e3: out <= 12'h000;
      20'h021e4: out <= 12'h000;
      20'h021e5: out <= 12'h000;
      20'h021e6: out <= 12'h000;
      20'h021e7: out <= 12'h000;
      20'h021e8: out <= 12'h000;
      20'h021e9: out <= 12'h000;
      20'h021ea: out <= 12'h000;
      20'h021eb: out <= 12'h000;
      20'h021ec: out <= 12'h000;
      20'h021ed: out <= 12'h000;
      20'h021ee: out <= 12'h000;
      20'h021ef: out <= 12'h000;
      20'h021f0: out <= 12'h000;
      20'h021f1: out <= 12'h000;
      20'h021f2: out <= 12'h000;
      20'h021f3: out <= 12'h000;
      20'h021f4: out <= 12'h000;
      20'h021f5: out <= 12'h000;
      20'h021f6: out <= 12'h000;
      20'h021f7: out <= 12'h000;
      20'h021f8: out <= 12'h222;
      20'h021f9: out <= 12'h222;
      20'h021fa: out <= 12'h222;
      20'h021fb: out <= 12'h222;
      20'h021fc: out <= 12'h222;
      20'h021fd: out <= 12'h222;
      20'h021fe: out <= 12'h222;
      20'h021ff: out <= 12'h222;
      20'h02200: out <= 12'h222;
      20'h02201: out <= 12'h222;
      20'h02202: out <= 12'h222;
      20'h02203: out <= 12'h222;
      20'h02204: out <= 12'h222;
      20'h02205: out <= 12'h222;
      20'h02206: out <= 12'h222;
      20'h02207: out <= 12'h222;
      20'h02208: out <= 12'h000;
      20'h02209: out <= 12'h000;
      20'h0220a: out <= 12'h000;
      20'h0220b: out <= 12'h000;
      20'h0220c: out <= 12'h000;
      20'h0220d: out <= 12'h000;
      20'h0220e: out <= 12'hfff;
      20'h0220f: out <= 12'hfff;
      20'h02210: out <= 12'hfff;
      20'h02211: out <= 12'hfff;
      20'h02212: out <= 12'hfff;
      20'h02213: out <= 12'h000;
      20'h02214: out <= 12'h000;
      20'h02215: out <= 12'h000;
      20'h02216: out <= 12'h000;
      20'h02217: out <= 12'h000;
      20'h02218: out <= 12'h222;
      20'h02219: out <= 12'h222;
      20'h0221a: out <= 12'h222;
      20'h0221b: out <= 12'h222;
      20'h0221c: out <= 12'h222;
      20'h0221d: out <= 12'h222;
      20'h0221e: out <= 12'h16d;
      20'h0221f: out <= 12'h16d;
      20'h02220: out <= 12'h16d;
      20'h02221: out <= 12'h16d;
      20'h02222: out <= 12'h16d;
      20'h02223: out <= 12'h222;
      20'h02224: out <= 12'h222;
      20'h02225: out <= 12'h222;
      20'h02226: out <= 12'h222;
      20'h02227: out <= 12'h222;
      20'h02228: out <= 12'h000;
      20'h02229: out <= 12'h000;
      20'h0222a: out <= 12'h000;
      20'h0222b: out <= 12'h000;
      20'h0222c: out <= 12'h000;
      20'h0222d: out <= 12'h000;
      20'h0222e: out <= 12'h000;
      20'h0222f: out <= 12'h000;
      20'h02230: out <= 12'h000;
      20'h02231: out <= 12'h000;
      20'h02232: out <= 12'h000;
      20'h02233: out <= 12'h000;
      20'h02234: out <= 12'h000;
      20'h02235: out <= 12'h000;
      20'h02236: out <= 12'h000;
      20'h02237: out <= 12'h000;
      20'h02238: out <= 12'h222;
      20'h02239: out <= 12'h222;
      20'h0223a: out <= 12'h222;
      20'h0223b: out <= 12'h222;
      20'h0223c: out <= 12'h222;
      20'h0223d: out <= 12'h222;
      20'h0223e: out <= 12'h222;
      20'h0223f: out <= 12'h222;
      20'h02240: out <= 12'h222;
      20'h02241: out <= 12'h222;
      20'h02242: out <= 12'h222;
      20'h02243: out <= 12'h222;
      20'h02244: out <= 12'h222;
      20'h02245: out <= 12'h222;
      20'h02246: out <= 12'h222;
      20'h02247: out <= 12'h222;
      20'h02248: out <= 12'h000;
      20'h02249: out <= 12'h000;
      20'h0224a: out <= 12'h000;
      20'h0224b: out <= 12'h000;
      20'h0224c: out <= 12'h000;
      20'h0224d: out <= 12'h000;
      20'h0224e: out <= 12'h000;
      20'h0224f: out <= 12'h6af;
      20'h02250: out <= 12'hfff;
      20'h02251: out <= 12'h6af;
      20'h02252: out <= 12'h000;
      20'h02253: out <= 12'h000;
      20'h02254: out <= 12'h000;
      20'h02255: out <= 12'h000;
      20'h02256: out <= 12'h000;
      20'h02257: out <= 12'h000;
      20'h02258: out <= 12'h222;
      20'h02259: out <= 12'h222;
      20'h0225a: out <= 12'h222;
      20'h0225b: out <= 12'h222;
      20'h0225c: out <= 12'h222;
      20'h0225d: out <= 12'h222;
      20'h0225e: out <= 12'h222;
      20'h0225f: out <= 12'h6af;
      20'h02260: out <= 12'hfff;
      20'h02261: out <= 12'h6af;
      20'h02262: out <= 12'h222;
      20'h02263: out <= 12'h222;
      20'h02264: out <= 12'h222;
      20'h02265: out <= 12'h222;
      20'h02266: out <= 12'h222;
      20'h02267: out <= 12'h222;
      20'h02268: out <= 12'h603;
      20'h02269: out <= 12'h603;
      20'h0226a: out <= 12'h603;
      20'h0226b: out <= 12'h603;
      20'h0226c: out <= 12'h666;
      20'h0226d: out <= 12'h666;
      20'h0226e: out <= 12'h666;
      20'h0226f: out <= 12'h666;
      20'h02270: out <= 12'h666;
      20'h02271: out <= 12'h666;
      20'h02272: out <= 12'h666;
      20'h02273: out <= 12'h666;
      20'h02274: out <= 12'h666;
      20'h02275: out <= 12'h666;
      20'h02276: out <= 12'h666;
      20'h02277: out <= 12'h666;
      20'h02278: out <= 12'h666;
      20'h02279: out <= 12'h666;
      20'h0227a: out <= 12'h666;
      20'h0227b: out <= 12'h666;
      20'h0227c: out <= 12'h000;
      20'h0227d: out <= 12'h000;
      20'h0227e: out <= 12'h000;
      20'h0227f: out <= 12'h000;
      20'h02280: out <= 12'h000;
      20'h02281: out <= 12'h000;
      20'h02282: out <= 12'h000;
      20'h02283: out <= 12'h000;
      20'h02284: out <= 12'h666;
      20'h02285: out <= 12'h666;
      20'h02286: out <= 12'h666;
      20'h02287: out <= 12'h666;
      20'h02288: out <= 12'h666;
      20'h02289: out <= 12'h666;
      20'h0228a: out <= 12'h666;
      20'h0228b: out <= 12'h666;
      20'h0228c: out <= 12'h666;
      20'h0228d: out <= 12'h666;
      20'h0228e: out <= 12'h666;
      20'h0228f: out <= 12'h666;
      20'h02290: out <= 12'h666;
      20'h02291: out <= 12'h666;
      20'h02292: out <= 12'h666;
      20'h02293: out <= 12'h666;
      20'h02294: out <= 12'h666;
      20'h02295: out <= 12'h666;
      20'h02296: out <= 12'h666;
      20'h02297: out <= 12'h666;
      20'h02298: out <= 12'h666;
      20'h02299: out <= 12'h666;
      20'h0229a: out <= 12'h666;
      20'h0229b: out <= 12'h666;
      20'h0229c: out <= 12'h666;
      20'h0229d: out <= 12'h666;
      20'h0229e: out <= 12'h666;
      20'h0229f: out <= 12'h666;
      20'h022a0: out <= 12'h666;
      20'h022a1: out <= 12'h666;
      20'h022a2: out <= 12'h666;
      20'h022a3: out <= 12'h666;
      20'h022a4: out <= 12'h000;
      20'h022a5: out <= 12'h000;
      20'h022a6: out <= 12'h000;
      20'h022a7: out <= 12'h000;
      20'h022a8: out <= 12'h000;
      20'h022a9: out <= 12'h000;
      20'h022aa: out <= 12'h000;
      20'h022ab: out <= 12'h000;
      20'h022ac: out <= 12'h000;
      20'h022ad: out <= 12'h000;
      20'h022ae: out <= 12'h000;
      20'h022af: out <= 12'h000;
      20'h022b0: out <= 12'h000;
      20'h022b1: out <= 12'h000;
      20'h022b2: out <= 12'h000;
      20'h022b3: out <= 12'h000;
      20'h022b4: out <= 12'h000;
      20'h022b5: out <= 12'h000;
      20'h022b6: out <= 12'h000;
      20'h022b7: out <= 12'h000;
      20'h022b8: out <= 12'h000;
      20'h022b9: out <= 12'h000;
      20'h022ba: out <= 12'h000;
      20'h022bb: out <= 12'h000;
      20'h022bc: out <= 12'h603;
      20'h022bd: out <= 12'h603;
      20'h022be: out <= 12'h603;
      20'h022bf: out <= 12'h603;
      20'h022c0: out <= 12'hb27;
      20'h022c1: out <= 12'hb27;
      20'h022c2: out <= 12'hb27;
      20'h022c3: out <= 12'hb27;
      20'h022c4: out <= 12'hb27;
      20'h022c5: out <= 12'hb27;
      20'h022c6: out <= 12'hb27;
      20'h022c7: out <= 12'hb27;
      20'h022c8: out <= 12'h000;
      20'h022c9: out <= 12'h000;
      20'h022ca: out <= 12'h000;
      20'h022cb: out <= 12'h000;
      20'h022cc: out <= 12'h000;
      20'h022cd: out <= 12'h000;
      20'h022ce: out <= 12'h000;
      20'h022cf: out <= 12'h000;
      20'h022d0: out <= 12'h000;
      20'h022d1: out <= 12'h000;
      20'h022d2: out <= 12'h000;
      20'h022d3: out <= 12'h000;
      20'h022d4: out <= 12'h000;
      20'h022d5: out <= 12'h000;
      20'h022d6: out <= 12'h000;
      20'h022d7: out <= 12'h000;
      20'h022d8: out <= 12'h000;
      20'h022d9: out <= 12'h000;
      20'h022da: out <= 12'h000;
      20'h022db: out <= 12'h000;
      20'h022dc: out <= 12'h000;
      20'h022dd: out <= 12'h000;
      20'h022de: out <= 12'h000;
      20'h022df: out <= 12'h000;
      20'h022e0: out <= 12'h000;
      20'h022e1: out <= 12'h000;
      20'h022e2: out <= 12'h000;
      20'h022e3: out <= 12'h000;
      20'h022e4: out <= 12'h000;
      20'h022e5: out <= 12'h000;
      20'h022e6: out <= 12'h000;
      20'h022e7: out <= 12'h000;
      20'h022e8: out <= 12'h000;
      20'h022e9: out <= 12'h000;
      20'h022ea: out <= 12'h000;
      20'h022eb: out <= 12'h000;
      20'h022ec: out <= 12'h000;
      20'h022ed: out <= 12'h000;
      20'h022ee: out <= 12'h000;
      20'h022ef: out <= 12'h000;
      20'h022f0: out <= 12'h000;
      20'h022f1: out <= 12'h000;
      20'h022f2: out <= 12'h000;
      20'h022f3: out <= 12'h000;
      20'h022f4: out <= 12'h000;
      20'h022f5: out <= 12'h000;
      20'h022f6: out <= 12'h000;
      20'h022f7: out <= 12'h000;
      20'h022f8: out <= 12'h000;
      20'h022f9: out <= 12'h000;
      20'h022fa: out <= 12'h000;
      20'h022fb: out <= 12'h000;
      20'h022fc: out <= 12'h000;
      20'h022fd: out <= 12'h000;
      20'h022fe: out <= 12'h000;
      20'h022ff: out <= 12'h000;
      20'h02300: out <= 12'h222;
      20'h02301: out <= 12'hc7f;
      20'h02302: out <= 12'hc7f;
      20'h02303: out <= 12'hc7f;
      20'h02304: out <= 12'hc7f;
      20'h02305: out <= 12'hc7f;
      20'h02306: out <= 12'hc7f;
      20'h02307: out <= 12'hc7f;
      20'h02308: out <= 12'hc7f;
      20'h02309: out <= 12'hc7f;
      20'h0230a: out <= 12'hc7f;
      20'h0230b: out <= 12'hc7f;
      20'h0230c: out <= 12'hc7f;
      20'h0230d: out <= 12'h222;
      20'h0230e: out <= 12'h222;
      20'h0230f: out <= 12'h222;
      20'h02310: out <= 12'h000;
      20'h02311: out <= 12'hc7f;
      20'h02312: out <= 12'hc7f;
      20'h02313: out <= 12'hc7f;
      20'h02314: out <= 12'hc7f;
      20'h02315: out <= 12'hc7f;
      20'h02316: out <= 12'hc7f;
      20'h02317: out <= 12'hc7f;
      20'h02318: out <= 12'hc7f;
      20'h02319: out <= 12'hc7f;
      20'h0231a: out <= 12'hc7f;
      20'h0231b: out <= 12'hc7f;
      20'h0231c: out <= 12'hc7f;
      20'h0231d: out <= 12'h000;
      20'h0231e: out <= 12'h000;
      20'h0231f: out <= 12'h000;
      20'h02320: out <= 12'h222;
      20'h02321: out <= 12'h222;
      20'h02322: out <= 12'h222;
      20'h02323: out <= 12'h222;
      20'h02324: out <= 12'h222;
      20'h02325: out <= 12'h222;
      20'h02326: out <= 12'h222;
      20'h02327: out <= 12'hc7f;
      20'h02328: out <= 12'hfff;
      20'h02329: out <= 12'hc7f;
      20'h0232a: out <= 12'h222;
      20'h0232b: out <= 12'h222;
      20'h0232c: out <= 12'h222;
      20'h0232d: out <= 12'h222;
      20'h0232e: out <= 12'h222;
      20'h0232f: out <= 12'h222;
      20'h02330: out <= 12'h000;
      20'h02331: out <= 12'h000;
      20'h02332: out <= 12'h000;
      20'h02333: out <= 12'h000;
      20'h02334: out <= 12'h000;
      20'h02335: out <= 12'h000;
      20'h02336: out <= 12'h000;
      20'h02337: out <= 12'hc7f;
      20'h02338: out <= 12'hfff;
      20'h02339: out <= 12'hc7f;
      20'h0233a: out <= 12'h000;
      20'h0233b: out <= 12'h000;
      20'h0233c: out <= 12'h000;
      20'h0233d: out <= 12'h000;
      20'h0233e: out <= 12'h000;
      20'h0233f: out <= 12'h000;
      20'h02340: out <= 12'h222;
      20'h02341: out <= 12'h222;
      20'h02342: out <= 12'h222;
      20'h02343: out <= 12'hc7f;
      20'h02344: out <= 12'hc7f;
      20'h02345: out <= 12'hc7f;
      20'h02346: out <= 12'hc7f;
      20'h02347: out <= 12'hc7f;
      20'h02348: out <= 12'hc7f;
      20'h02349: out <= 12'hc7f;
      20'h0234a: out <= 12'hc7f;
      20'h0234b: out <= 12'hc7f;
      20'h0234c: out <= 12'hc7f;
      20'h0234d: out <= 12'hc7f;
      20'h0234e: out <= 12'hc7f;
      20'h0234f: out <= 12'h222;
      20'h02350: out <= 12'h000;
      20'h02351: out <= 12'h000;
      20'h02352: out <= 12'h000;
      20'h02353: out <= 12'hc7f;
      20'h02354: out <= 12'hc7f;
      20'h02355: out <= 12'hc7f;
      20'h02356: out <= 12'hc7f;
      20'h02357: out <= 12'hc7f;
      20'h02358: out <= 12'hc7f;
      20'h02359: out <= 12'hc7f;
      20'h0235a: out <= 12'hc7f;
      20'h0235b: out <= 12'hc7f;
      20'h0235c: out <= 12'hc7f;
      20'h0235d: out <= 12'hc7f;
      20'h0235e: out <= 12'hc7f;
      20'h0235f: out <= 12'h000;
      20'h02360: out <= 12'h222;
      20'h02361: out <= 12'h222;
      20'h02362: out <= 12'h222;
      20'h02363: out <= 12'h222;
      20'h02364: out <= 12'h222;
      20'h02365: out <= 12'h222;
      20'h02366: out <= 12'h222;
      20'h02367: out <= 12'h222;
      20'h02368: out <= 12'h222;
      20'h02369: out <= 12'h222;
      20'h0236a: out <= 12'h222;
      20'h0236b: out <= 12'h222;
      20'h0236c: out <= 12'h222;
      20'h0236d: out <= 12'h222;
      20'h0236e: out <= 12'h222;
      20'h0236f: out <= 12'h222;
      20'h02370: out <= 12'h000;
      20'h02371: out <= 12'h000;
      20'h02372: out <= 12'h000;
      20'h02373: out <= 12'h000;
      20'h02374: out <= 12'h000;
      20'h02375: out <= 12'h000;
      20'h02376: out <= 12'h000;
      20'h02377: out <= 12'h000;
      20'h02378: out <= 12'h000;
      20'h02379: out <= 12'h000;
      20'h0237a: out <= 12'h000;
      20'h0237b: out <= 12'h000;
      20'h0237c: out <= 12'h000;
      20'h0237d: out <= 12'h000;
      20'h0237e: out <= 12'h000;
      20'h0237f: out <= 12'h000;
      20'h02380: out <= 12'h603;
      20'h02381: out <= 12'h603;
      20'h02382: out <= 12'h603;
      20'h02383: out <= 12'h603;
      20'h02384: out <= 12'hfff;
      20'h02385: out <= 12'h6af;
      20'h02386: out <= 12'h6af;
      20'h02387: out <= 12'hfff;
      20'h02388: out <= 12'h4cd;
      20'h02389: out <= 12'h4cd;
      20'h0238a: out <= 12'h4cd;
      20'h0238b: out <= 12'h4cd;
      20'h0238c: out <= 12'hfff;
      20'h0238d: out <= 12'h6af;
      20'h0238e: out <= 12'h6af;
      20'h0238f: out <= 12'hfff;
      20'h02390: out <= 12'h4cd;
      20'h02391: out <= 12'h4cd;
      20'h02392: out <= 12'h4cd;
      20'h02393: out <= 12'h4cd;
      20'h02394: out <= 12'h000;
      20'h02395: out <= 12'h000;
      20'h02396: out <= 12'hfff;
      20'h02397: out <= 12'hfff;
      20'h02398: out <= 12'hfff;
      20'h02399: out <= 12'h8d0;
      20'h0239a: out <= 12'h380;
      20'h0239b: out <= 12'h000;
      20'h0239c: out <= 12'h000;
      20'h0239d: out <= 12'h000;
      20'h0239e: out <= 12'hfff;
      20'h0239f: out <= 12'hfff;
      20'h023a0: out <= 12'hfff;
      20'h023a1: out <= 12'h8d0;
      20'h023a2: out <= 12'h380;
      20'h023a3: out <= 12'h000;
      20'h023a4: out <= 12'hfff;
      20'h023a5: out <= 12'h666;
      20'h023a6: out <= 12'h000;
      20'h023a7: out <= 12'h000;
      20'h023a8: out <= 12'hfff;
      20'h023a9: out <= 12'h666;
      20'h023aa: out <= 12'h000;
      20'h023ab: out <= 12'h000;
      20'h023ac: out <= 12'hfff;
      20'h023ad: out <= 12'h666;
      20'h023ae: out <= 12'h000;
      20'h023af: out <= 12'h000;
      20'h023b0: out <= 12'hfff;
      20'h023b1: out <= 12'h666;
      20'h023b2: out <= 12'h000;
      20'h023b3: out <= 12'h000;
      20'h023b4: out <= 12'h000;
      20'h023b5: out <= 12'h000;
      20'h023b6: out <= 12'h000;
      20'h023b7: out <= 12'h000;
      20'h023b8: out <= 12'h000;
      20'h023b9: out <= 12'h000;
      20'h023ba: out <= 12'h000;
      20'h023bb: out <= 12'h000;
      20'h023bc: out <= 12'h6af;
      20'h023bd: out <= 12'h6af;
      20'h023be: out <= 12'h000;
      20'h023bf: out <= 12'h000;
      20'h023c0: out <= 12'h000;
      20'h023c1: out <= 12'h000;
      20'h023c2: out <= 12'h000;
      20'h023c3: out <= 12'h000;
      20'h023c4: out <= 12'h000;
      20'h023c5: out <= 12'h000;
      20'h023c6: out <= 12'h000;
      20'h023c7: out <= 12'h000;
      20'h023c8: out <= 12'h000;
      20'h023c9: out <= 12'h000;
      20'h023ca: out <= 12'h000;
      20'h023cb: out <= 12'h000;
      20'h023cc: out <= 12'h000;
      20'h023cd: out <= 12'h000;
      20'h023ce: out <= 12'h000;
      20'h023cf: out <= 12'h000;
      20'h023d0: out <= 12'h000;
      20'h023d1: out <= 12'h000;
      20'h023d2: out <= 12'h000;
      20'h023d3: out <= 12'h000;
      20'h023d4: out <= 12'h603;
      20'h023d5: out <= 12'h603;
      20'h023d6: out <= 12'h603;
      20'h023d7: out <= 12'h603;
      20'h023d8: out <= 12'hee9;
      20'h023d9: out <= 12'hee9;
      20'h023da: out <= 12'hee9;
      20'h023db: out <= 12'hee9;
      20'h023dc: out <= 12'hee9;
      20'h023dd: out <= 12'hee9;
      20'h023de: out <= 12'hee9;
      20'h023df: out <= 12'hb27;
      20'h023e0: out <= 12'h000;
      20'h023e1: out <= 12'h000;
      20'h023e2: out <= 12'h000;
      20'h023e3: out <= 12'h000;
      20'h023e4: out <= 12'h000;
      20'h023e5: out <= 12'h000;
      20'h023e6: out <= 12'h000;
      20'h023e7: out <= 12'h000;
      20'h023e8: out <= 12'h000;
      20'h023e9: out <= 12'h000;
      20'h023ea: out <= 12'h000;
      20'h023eb: out <= 12'h000;
      20'h023ec: out <= 12'h000;
      20'h023ed: out <= 12'h000;
      20'h023ee: out <= 12'h000;
      20'h023ef: out <= 12'h000;
      20'h023f0: out <= 12'h916;
      20'h023f1: out <= 12'h916;
      20'h023f2: out <= 12'h916;
      20'h023f3: out <= 12'h916;
      20'h023f4: out <= 12'h916;
      20'h023f5: out <= 12'h916;
      20'h023f6: out <= 12'h916;
      20'h023f7: out <= 12'h916;
      20'h023f8: out <= 12'hd29;
      20'h023f9: out <= 12'hd29;
      20'h023fa: out <= 12'hd29;
      20'h023fb: out <= 12'hd29;
      20'h023fc: out <= 12'hd29;
      20'h023fd: out <= 12'hd29;
      20'h023fe: out <= 12'hd29;
      20'h023ff: out <= 12'hd29;
      20'h02400: out <= 12'h000;
      20'h02401: out <= 12'h000;
      20'h02402: out <= 12'h000;
      20'h02403: out <= 12'h000;
      20'h02404: out <= 12'h000;
      20'h02405: out <= 12'h000;
      20'h02406: out <= 12'h000;
      20'h02407: out <= 12'h000;
      20'h02408: out <= 12'h000;
      20'h02409: out <= 12'h000;
      20'h0240a: out <= 12'h000;
      20'h0240b: out <= 12'h000;
      20'h0240c: out <= 12'h000;
      20'h0240d: out <= 12'h000;
      20'h0240e: out <= 12'h000;
      20'h0240f: out <= 12'h000;
      20'h02410: out <= 12'h000;
      20'h02411: out <= 12'h000;
      20'h02412: out <= 12'h000;
      20'h02413: out <= 12'h000;
      20'h02414: out <= 12'h000;
      20'h02415: out <= 12'h000;
      20'h02416: out <= 12'h000;
      20'h02417: out <= 12'h000;
      20'h02418: out <= 12'h222;
      20'h02419: out <= 12'hfff;
      20'h0241a: out <= 12'h72f;
      20'h0241b: out <= 12'hfff;
      20'h0241c: out <= 12'h72f;
      20'h0241d: out <= 12'hfff;
      20'h0241e: out <= 12'h72f;
      20'h0241f: out <= 12'hfff;
      20'h02420: out <= 12'h72f;
      20'h02421: out <= 12'hfff;
      20'h02422: out <= 12'h72f;
      20'h02423: out <= 12'hfff;
      20'h02424: out <= 12'h72f;
      20'h02425: out <= 12'h222;
      20'h02426: out <= 12'h222;
      20'h02427: out <= 12'h222;
      20'h02428: out <= 12'h000;
      20'h02429: out <= 12'hc7f;
      20'h0242a: out <= 12'hfff;
      20'h0242b: out <= 12'h72f;
      20'h0242c: out <= 12'hfff;
      20'h0242d: out <= 12'h72f;
      20'h0242e: out <= 12'hfff;
      20'h0242f: out <= 12'h72f;
      20'h02430: out <= 12'hfff;
      20'h02431: out <= 12'h72f;
      20'h02432: out <= 12'hfff;
      20'h02433: out <= 12'h72f;
      20'h02434: out <= 12'hfff;
      20'h02435: out <= 12'h000;
      20'h02436: out <= 12'h000;
      20'h02437: out <= 12'h000;
      20'h02438: out <= 12'h222;
      20'h02439: out <= 12'h222;
      20'h0243a: out <= 12'h222;
      20'h0243b: out <= 12'h222;
      20'h0243c: out <= 12'h222;
      20'h0243d: out <= 12'h222;
      20'h0243e: out <= 12'h222;
      20'h0243f: out <= 12'h72f;
      20'h02440: out <= 12'hfff;
      20'h02441: out <= 12'h72f;
      20'h02442: out <= 12'h222;
      20'h02443: out <= 12'h222;
      20'h02444: out <= 12'h222;
      20'h02445: out <= 12'h222;
      20'h02446: out <= 12'h222;
      20'h02447: out <= 12'h222;
      20'h02448: out <= 12'h000;
      20'h02449: out <= 12'h000;
      20'h0244a: out <= 12'h000;
      20'h0244b: out <= 12'h000;
      20'h0244c: out <= 12'h000;
      20'h0244d: out <= 12'h000;
      20'h0244e: out <= 12'h000;
      20'h0244f: out <= 12'h72f;
      20'h02450: out <= 12'hfff;
      20'h02451: out <= 12'h72f;
      20'h02452: out <= 12'h000;
      20'h02453: out <= 12'h000;
      20'h02454: out <= 12'h000;
      20'h02455: out <= 12'h000;
      20'h02456: out <= 12'h000;
      20'h02457: out <= 12'h000;
      20'h02458: out <= 12'h222;
      20'h02459: out <= 12'h222;
      20'h0245a: out <= 12'h222;
      20'h0245b: out <= 12'h72f;
      20'h0245c: out <= 12'hfff;
      20'h0245d: out <= 12'h72f;
      20'h0245e: out <= 12'hfff;
      20'h0245f: out <= 12'h72f;
      20'h02460: out <= 12'hfff;
      20'h02461: out <= 12'h72f;
      20'h02462: out <= 12'hfff;
      20'h02463: out <= 12'h72f;
      20'h02464: out <= 12'hfff;
      20'h02465: out <= 12'h72f;
      20'h02466: out <= 12'hfff;
      20'h02467: out <= 12'h222;
      20'h02468: out <= 12'h000;
      20'h02469: out <= 12'h000;
      20'h0246a: out <= 12'h000;
      20'h0246b: out <= 12'hfff;
      20'h0246c: out <= 12'h72f;
      20'h0246d: out <= 12'hfff;
      20'h0246e: out <= 12'h72f;
      20'h0246f: out <= 12'hfff;
      20'h02470: out <= 12'h72f;
      20'h02471: out <= 12'hfff;
      20'h02472: out <= 12'h72f;
      20'h02473: out <= 12'hfff;
      20'h02474: out <= 12'h72f;
      20'h02475: out <= 12'hfff;
      20'h02476: out <= 12'hc7f;
      20'h02477: out <= 12'h000;
      20'h02478: out <= 12'h222;
      20'h02479: out <= 12'hc7f;
      20'h0247a: out <= 12'hfff;
      20'h0247b: out <= 12'hc7f;
      20'h0247c: out <= 12'h222;
      20'h0247d: out <= 12'h222;
      20'h0247e: out <= 12'h222;
      20'h0247f: out <= 12'h222;
      20'h02480: out <= 12'h222;
      20'h02481: out <= 12'h222;
      20'h02482: out <= 12'h222;
      20'h02483: out <= 12'h222;
      20'h02484: out <= 12'h222;
      20'h02485: out <= 12'hc7f;
      20'h02486: out <= 12'hfff;
      20'h02487: out <= 12'hc7f;
      20'h02488: out <= 12'h000;
      20'h02489: out <= 12'hc7f;
      20'h0248a: out <= 12'hc7f;
      20'h0248b: out <= 12'hc7f;
      20'h0248c: out <= 12'h000;
      20'h0248d: out <= 12'h000;
      20'h0248e: out <= 12'h000;
      20'h0248f: out <= 12'h000;
      20'h02490: out <= 12'h000;
      20'h02491: out <= 12'h000;
      20'h02492: out <= 12'h000;
      20'h02493: out <= 12'h000;
      20'h02494: out <= 12'h000;
      20'h02495: out <= 12'hc7f;
      20'h02496: out <= 12'hc7f;
      20'h02497: out <= 12'hc7f;
      20'h02498: out <= 12'h603;
      20'h02499: out <= 12'h603;
      20'h0249a: out <= 12'h603;
      20'h0249b: out <= 12'h603;
      20'h0249c: out <= 12'h4cd;
      20'h0249d: out <= 12'hfff;
      20'h0249e: out <= 12'hfff;
      20'h0249f: out <= 12'h4cd;
      20'h024a0: out <= 12'h4cd;
      20'h024a1: out <= 12'h6af;
      20'h024a2: out <= 12'h6af;
      20'h024a3: out <= 12'h4cd;
      20'h024a4: out <= 12'h4cd;
      20'h024a5: out <= 12'hfff;
      20'h024a6: out <= 12'hfff;
      20'h024a7: out <= 12'h4cd;
      20'h024a8: out <= 12'h4cd;
      20'h024a9: out <= 12'h6af;
      20'h024aa: out <= 12'h6af;
      20'h024ab: out <= 12'h4cd;
      20'h024ac: out <= 12'h000;
      20'h024ad: out <= 12'hfff;
      20'h024ae: out <= 12'h8d0;
      20'h024af: out <= 12'hfff;
      20'h024b0: out <= 12'h8d0;
      20'h024b1: out <= 12'h380;
      20'h024b2: out <= 12'h8d0;
      20'h024b3: out <= 12'h380;
      20'h024b4: out <= 12'h000;
      20'h024b5: out <= 12'hfff;
      20'h024b6: out <= 12'h8d0;
      20'h024b7: out <= 12'hfff;
      20'h024b8: out <= 12'h8d0;
      20'h024b9: out <= 12'h380;
      20'h024ba: out <= 12'h8d0;
      20'h024bb: out <= 12'h380;
      20'h024bc: out <= 12'hbbb;
      20'h024bd: out <= 12'hfff;
      20'h024be: out <= 12'h000;
      20'h024bf: out <= 12'h000;
      20'h024c0: out <= 12'hbbb;
      20'h024c1: out <= 12'hfff;
      20'h024c2: out <= 12'h000;
      20'h024c3: out <= 12'h000;
      20'h024c4: out <= 12'hbbb;
      20'h024c5: out <= 12'hfff;
      20'h024c6: out <= 12'h000;
      20'h024c7: out <= 12'h000;
      20'h024c8: out <= 12'hbbb;
      20'h024c9: out <= 12'hfff;
      20'h024ca: out <= 12'h000;
      20'h024cb: out <= 12'h000;
      20'h024cc: out <= 12'h000;
      20'h024cd: out <= 12'h000;
      20'h024ce: out <= 12'h000;
      20'h024cf: out <= 12'h000;
      20'h024d0: out <= 12'h000;
      20'h024d1: out <= 12'h000;
      20'h024d2: out <= 12'h000;
      20'h024d3: out <= 12'h6af;
      20'h024d4: out <= 12'h4cd;
      20'h024d5: out <= 12'h4cd;
      20'h024d6: out <= 12'h6af;
      20'h024d7: out <= 12'h000;
      20'h024d8: out <= 12'h000;
      20'h024d9: out <= 12'h000;
      20'h024da: out <= 12'h000;
      20'h024db: out <= 12'h000;
      20'h024dc: out <= 12'h000;
      20'h024dd: out <= 12'h000;
      20'h024de: out <= 12'h000;
      20'h024df: out <= 12'h000;
      20'h024e0: out <= 12'h000;
      20'h024e1: out <= 12'h000;
      20'h024e2: out <= 12'h000;
      20'h024e3: out <= 12'h000;
      20'h024e4: out <= 12'h000;
      20'h024e5: out <= 12'h000;
      20'h024e6: out <= 12'h000;
      20'h024e7: out <= 12'h000;
      20'h024e8: out <= 12'h000;
      20'h024e9: out <= 12'h000;
      20'h024ea: out <= 12'h000;
      20'h024eb: out <= 12'h000;
      20'h024ec: out <= 12'h603;
      20'h024ed: out <= 12'h603;
      20'h024ee: out <= 12'h603;
      20'h024ef: out <= 12'h603;
      20'h024f0: out <= 12'hee9;
      20'h024f1: out <= 12'hf87;
      20'h024f2: out <= 12'hf87;
      20'h024f3: out <= 12'hf87;
      20'h024f4: out <= 12'hf87;
      20'h024f5: out <= 12'hf87;
      20'h024f6: out <= 12'hf87;
      20'h024f7: out <= 12'hb27;
      20'h024f8: out <= 12'h000;
      20'h024f9: out <= 12'h000;
      20'h024fa: out <= 12'h000;
      20'h024fb: out <= 12'h000;
      20'h024fc: out <= 12'h000;
      20'h024fd: out <= 12'h000;
      20'h024fe: out <= 12'h000;
      20'h024ff: out <= 12'h000;
      20'h02500: out <= 12'h000;
      20'h02501: out <= 12'h000;
      20'h02502: out <= 12'h000;
      20'h02503: out <= 12'h000;
      20'h02504: out <= 12'h000;
      20'h02505: out <= 12'h000;
      20'h02506: out <= 12'h000;
      20'h02507: out <= 12'h000;
      20'h02508: out <= 12'h916;
      20'h02509: out <= 12'h916;
      20'h0250a: out <= 12'h916;
      20'h0250b: out <= 12'h916;
      20'h0250c: out <= 12'h916;
      20'h0250d: out <= 12'h916;
      20'h0250e: out <= 12'h916;
      20'h0250f: out <= 12'h916;
      20'h02510: out <= 12'hd29;
      20'h02511: out <= 12'hd29;
      20'h02512: out <= 12'hd29;
      20'h02513: out <= 12'hd29;
      20'h02514: out <= 12'hd29;
      20'h02515: out <= 12'hd29;
      20'h02516: out <= 12'hd29;
      20'h02517: out <= 12'hd29;
      20'h02518: out <= 12'h000;
      20'h02519: out <= 12'h000;
      20'h0251a: out <= 12'h000;
      20'h0251b: out <= 12'h000;
      20'h0251c: out <= 12'h000;
      20'h0251d: out <= 12'h000;
      20'h0251e: out <= 12'h000;
      20'h0251f: out <= 12'h000;
      20'h02520: out <= 12'h000;
      20'h02521: out <= 12'h000;
      20'h02522: out <= 12'h000;
      20'h02523: out <= 12'h000;
      20'h02524: out <= 12'h000;
      20'h02525: out <= 12'h000;
      20'h02526: out <= 12'h000;
      20'h02527: out <= 12'h000;
      20'h02528: out <= 12'h000;
      20'h02529: out <= 12'h000;
      20'h0252a: out <= 12'h000;
      20'h0252b: out <= 12'h000;
      20'h0252c: out <= 12'h000;
      20'h0252d: out <= 12'h000;
      20'h0252e: out <= 12'h000;
      20'h0252f: out <= 12'h000;
      20'h02530: out <= 12'h222;
      20'h02531: out <= 12'hc7f;
      20'h02532: out <= 12'hc7f;
      20'h02533: out <= 12'hc7f;
      20'h02534: out <= 12'h72f;
      20'h02535: out <= 12'h72f;
      20'h02536: out <= 12'h72f;
      20'h02537: out <= 12'h72f;
      20'h02538: out <= 12'h72f;
      20'h02539: out <= 12'h72f;
      20'h0253a: out <= 12'h72f;
      20'h0253b: out <= 12'hc7f;
      20'h0253c: out <= 12'hc7f;
      20'h0253d: out <= 12'h222;
      20'h0253e: out <= 12'h222;
      20'h0253f: out <= 12'h222;
      20'h02540: out <= 12'h000;
      20'h02541: out <= 12'hc7f;
      20'h02542: out <= 12'hc7f;
      20'h02543: out <= 12'hc7f;
      20'h02544: out <= 12'h72f;
      20'h02545: out <= 12'h72f;
      20'h02546: out <= 12'h72f;
      20'h02547: out <= 12'h72f;
      20'h02548: out <= 12'h72f;
      20'h02549: out <= 12'h72f;
      20'h0254a: out <= 12'h72f;
      20'h0254b: out <= 12'hc7f;
      20'h0254c: out <= 12'hc7f;
      20'h0254d: out <= 12'h000;
      20'h0254e: out <= 12'h000;
      20'h0254f: out <= 12'h000;
      20'h02550: out <= 12'h222;
      20'h02551: out <= 12'h222;
      20'h02552: out <= 12'h222;
      20'h02553: out <= 12'h222;
      20'h02554: out <= 12'h222;
      20'h02555: out <= 12'h222;
      20'h02556: out <= 12'h222;
      20'h02557: out <= 12'h72f;
      20'h02558: out <= 12'hfff;
      20'h02559: out <= 12'h72f;
      20'h0255a: out <= 12'h222;
      20'h0255b: out <= 12'h222;
      20'h0255c: out <= 12'h222;
      20'h0255d: out <= 12'h222;
      20'h0255e: out <= 12'h222;
      20'h0255f: out <= 12'h222;
      20'h02560: out <= 12'h000;
      20'h02561: out <= 12'h000;
      20'h02562: out <= 12'h000;
      20'h02563: out <= 12'h000;
      20'h02564: out <= 12'h000;
      20'h02565: out <= 12'h000;
      20'h02566: out <= 12'h000;
      20'h02567: out <= 12'h72f;
      20'h02568: out <= 12'hfff;
      20'h02569: out <= 12'h72f;
      20'h0256a: out <= 12'h000;
      20'h0256b: out <= 12'h000;
      20'h0256c: out <= 12'h000;
      20'h0256d: out <= 12'h000;
      20'h0256e: out <= 12'h000;
      20'h0256f: out <= 12'h000;
      20'h02570: out <= 12'h222;
      20'h02571: out <= 12'h222;
      20'h02572: out <= 12'h222;
      20'h02573: out <= 12'hc7f;
      20'h02574: out <= 12'hc7f;
      20'h02575: out <= 12'h72f;
      20'h02576: out <= 12'h72f;
      20'h02577: out <= 12'h72f;
      20'h02578: out <= 12'h72f;
      20'h02579: out <= 12'h72f;
      20'h0257a: out <= 12'h72f;
      20'h0257b: out <= 12'h72f;
      20'h0257c: out <= 12'hc7f;
      20'h0257d: out <= 12'hc7f;
      20'h0257e: out <= 12'hc7f;
      20'h0257f: out <= 12'h222;
      20'h02580: out <= 12'h000;
      20'h02581: out <= 12'h000;
      20'h02582: out <= 12'h000;
      20'h02583: out <= 12'hc7f;
      20'h02584: out <= 12'hc7f;
      20'h02585: out <= 12'h72f;
      20'h02586: out <= 12'h72f;
      20'h02587: out <= 12'h72f;
      20'h02588: out <= 12'h72f;
      20'h02589: out <= 12'h72f;
      20'h0258a: out <= 12'h72f;
      20'h0258b: out <= 12'h72f;
      20'h0258c: out <= 12'hc7f;
      20'h0258d: out <= 12'hc7f;
      20'h0258e: out <= 12'hc7f;
      20'h0258f: out <= 12'h000;
      20'h02590: out <= 12'h222;
      20'h02591: out <= 12'hc7f;
      20'h02592: out <= 12'h72f;
      20'h02593: out <= 12'hc7f;
      20'h02594: out <= 12'h222;
      20'h02595: out <= 12'h72f;
      20'h02596: out <= 12'h72f;
      20'h02597: out <= 12'h72f;
      20'h02598: out <= 12'h72f;
      20'h02599: out <= 12'h72f;
      20'h0259a: out <= 12'h72f;
      20'h0259b: out <= 12'h72f;
      20'h0259c: out <= 12'h222;
      20'h0259d: out <= 12'hc7f;
      20'h0259e: out <= 12'h72f;
      20'h0259f: out <= 12'hc7f;
      20'h025a0: out <= 12'h000;
      20'h025a1: out <= 12'hc7f;
      20'h025a2: out <= 12'hfff;
      20'h025a3: out <= 12'hc7f;
      20'h025a4: out <= 12'h000;
      20'h025a5: out <= 12'h72f;
      20'h025a6: out <= 12'h72f;
      20'h025a7: out <= 12'h72f;
      20'h025a8: out <= 12'h72f;
      20'h025a9: out <= 12'h72f;
      20'h025aa: out <= 12'h72f;
      20'h025ab: out <= 12'h72f;
      20'h025ac: out <= 12'h000;
      20'h025ad: out <= 12'hc7f;
      20'h025ae: out <= 12'hfff;
      20'h025af: out <= 12'hc7f;
      20'h025b0: out <= 12'h603;
      20'h025b1: out <= 12'h603;
      20'h025b2: out <= 12'h603;
      20'h025b3: out <= 12'h603;
      20'h025b4: out <= 12'h4cd;
      20'h025b5: out <= 12'h4cd;
      20'h025b6: out <= 12'h4cd;
      20'h025b7: out <= 12'h4cd;
      20'h025b8: out <= 12'h6af;
      20'h025b9: out <= 12'hfff;
      20'h025ba: out <= 12'hfff;
      20'h025bb: out <= 12'h6af;
      20'h025bc: out <= 12'h4cd;
      20'h025bd: out <= 12'h4cd;
      20'h025be: out <= 12'h4cd;
      20'h025bf: out <= 12'h4cd;
      20'h025c0: out <= 12'h6af;
      20'h025c1: out <= 12'hfff;
      20'h025c2: out <= 12'hfff;
      20'h025c3: out <= 12'h6af;
      20'h025c4: out <= 12'hfff;
      20'h025c5: out <= 12'h8d0;
      20'h025c6: out <= 12'hfff;
      20'h025c7: out <= 12'h8d0;
      20'h025c8: out <= 12'h8d0;
      20'h025c9: out <= 12'h8d0;
      20'h025ca: out <= 12'h380;
      20'h025cb: out <= 12'h8d0;
      20'h025cc: out <= 12'hfff;
      20'h025cd: out <= 12'h8d0;
      20'h025ce: out <= 12'hfff;
      20'h025cf: out <= 12'h8d0;
      20'h025d0: out <= 12'h8d0;
      20'h025d1: out <= 12'h8d0;
      20'h025d2: out <= 12'h380;
      20'h025d3: out <= 12'h8d0;
      20'h025d4: out <= 12'h000;
      20'h025d5: out <= 12'h000;
      20'h025d6: out <= 12'hfff;
      20'h025d7: out <= 12'h666;
      20'h025d8: out <= 12'h000;
      20'h025d9: out <= 12'h000;
      20'h025da: out <= 12'hfff;
      20'h025db: out <= 12'h666;
      20'h025dc: out <= 12'h000;
      20'h025dd: out <= 12'h000;
      20'h025de: out <= 12'hfff;
      20'h025df: out <= 12'h666;
      20'h025e0: out <= 12'h000;
      20'h025e1: out <= 12'h000;
      20'h025e2: out <= 12'hfff;
      20'h025e3: out <= 12'h666;
      20'h025e4: out <= 12'h000;
      20'h025e5: out <= 12'h000;
      20'h025e6: out <= 12'h000;
      20'h025e7: out <= 12'h000;
      20'h025e8: out <= 12'h000;
      20'h025e9: out <= 12'h000;
      20'h025ea: out <= 12'h6af;
      20'h025eb: out <= 12'h4cd;
      20'h025ec: out <= 12'hfff;
      20'h025ed: out <= 12'hfff;
      20'h025ee: out <= 12'h4cd;
      20'h025ef: out <= 12'h6af;
      20'h025f0: out <= 12'h000;
      20'h025f1: out <= 12'h000;
      20'h025f2: out <= 12'h000;
      20'h025f3: out <= 12'h000;
      20'h025f4: out <= 12'h000;
      20'h025f5: out <= 12'h000;
      20'h025f6: out <= 12'h000;
      20'h025f7: out <= 12'h000;
      20'h025f8: out <= 12'h000;
      20'h025f9: out <= 12'h000;
      20'h025fa: out <= 12'h000;
      20'h025fb: out <= 12'h000;
      20'h025fc: out <= 12'h000;
      20'h025fd: out <= 12'h000;
      20'h025fe: out <= 12'h6af;
      20'h025ff: out <= 12'h6af;
      20'h02600: out <= 12'h6af;
      20'h02601: out <= 12'h6af;
      20'h02602: out <= 12'h6af;
      20'h02603: out <= 12'h000;
      20'h02604: out <= 12'h603;
      20'h02605: out <= 12'h603;
      20'h02606: out <= 12'h603;
      20'h02607: out <= 12'h603;
      20'h02608: out <= 12'hee9;
      20'h02609: out <= 12'hf87;
      20'h0260a: out <= 12'hee9;
      20'h0260b: out <= 12'hee9;
      20'h0260c: out <= 12'hee9;
      20'h0260d: out <= 12'hb27;
      20'h0260e: out <= 12'hf87;
      20'h0260f: out <= 12'hb27;
      20'h02610: out <= 12'h000;
      20'h02611: out <= 12'h000;
      20'h02612: out <= 12'h000;
      20'h02613: out <= 12'h000;
      20'h02614: out <= 12'h000;
      20'h02615: out <= 12'h000;
      20'h02616: out <= 12'h000;
      20'h02617: out <= 12'h000;
      20'h02618: out <= 12'h000;
      20'h02619: out <= 12'h000;
      20'h0261a: out <= 12'h000;
      20'h0261b: out <= 12'h000;
      20'h0261c: out <= 12'h000;
      20'h0261d: out <= 12'h000;
      20'h0261e: out <= 12'h000;
      20'h0261f: out <= 12'h000;
      20'h02620: out <= 12'h916;
      20'h02621: out <= 12'h916;
      20'h02622: out <= 12'h916;
      20'h02623: out <= 12'h916;
      20'h02624: out <= 12'h916;
      20'h02625: out <= 12'h916;
      20'h02626: out <= 12'h916;
      20'h02627: out <= 12'h916;
      20'h02628: out <= 12'hd29;
      20'h02629: out <= 12'hd29;
      20'h0262a: out <= 12'hd29;
      20'h0262b: out <= 12'hd29;
      20'h0262c: out <= 12'hd29;
      20'h0262d: out <= 12'hd29;
      20'h0262e: out <= 12'hd29;
      20'h0262f: out <= 12'hd29;
      20'h02630: out <= 12'h000;
      20'h02631: out <= 12'h000;
      20'h02632: out <= 12'h000;
      20'h02633: out <= 12'h000;
      20'h02634: out <= 12'h000;
      20'h02635: out <= 12'h000;
      20'h02636: out <= 12'h000;
      20'h02637: out <= 12'h000;
      20'h02638: out <= 12'h000;
      20'h02639: out <= 12'h000;
      20'h0263a: out <= 12'h000;
      20'h0263b: out <= 12'h000;
      20'h0263c: out <= 12'h000;
      20'h0263d: out <= 12'h000;
      20'h0263e: out <= 12'h000;
      20'h0263f: out <= 12'h000;
      20'h02640: out <= 12'h000;
      20'h02641: out <= 12'h000;
      20'h02642: out <= 12'h000;
      20'h02643: out <= 12'h000;
      20'h02644: out <= 12'h000;
      20'h02645: out <= 12'h000;
      20'h02646: out <= 12'h000;
      20'h02647: out <= 12'h000;
      20'h02648: out <= 12'h222;
      20'h02649: out <= 12'h222;
      20'h0264a: out <= 12'h222;
      20'h0264b: out <= 12'h72f;
      20'h0264c: out <= 12'hfff;
      20'h0264d: out <= 12'hc7f;
      20'h0264e: out <= 12'hc7f;
      20'h0264f: out <= 12'hc7f;
      20'h02650: out <= 12'hc7f;
      20'h02651: out <= 12'hfff;
      20'h02652: out <= 12'h72f;
      20'h02653: out <= 12'h222;
      20'h02654: out <= 12'h222;
      20'h02655: out <= 12'h222;
      20'h02656: out <= 12'h222;
      20'h02657: out <= 12'h222;
      20'h02658: out <= 12'h000;
      20'h02659: out <= 12'h000;
      20'h0265a: out <= 12'h000;
      20'h0265b: out <= 12'h72f;
      20'h0265c: out <= 12'hfff;
      20'h0265d: out <= 12'hc7f;
      20'h0265e: out <= 12'hc7f;
      20'h0265f: out <= 12'hc7f;
      20'h02660: out <= 12'hc7f;
      20'h02661: out <= 12'hfff;
      20'h02662: out <= 12'h72f;
      20'h02663: out <= 12'h000;
      20'h02664: out <= 12'h000;
      20'h02665: out <= 12'h000;
      20'h02666: out <= 12'h000;
      20'h02667: out <= 12'h000;
      20'h02668: out <= 12'h222;
      20'h02669: out <= 12'hc7f;
      20'h0266a: out <= 12'h72f;
      20'h0266b: out <= 12'hc7f;
      20'h0266c: out <= 12'h222;
      20'h0266d: out <= 12'h222;
      20'h0266e: out <= 12'h222;
      20'h0266f: out <= 12'h72f;
      20'h02670: out <= 12'hfff;
      20'h02671: out <= 12'h72f;
      20'h02672: out <= 12'h222;
      20'h02673: out <= 12'h222;
      20'h02674: out <= 12'h222;
      20'h02675: out <= 12'hc7f;
      20'h02676: out <= 12'h72f;
      20'h02677: out <= 12'hc7f;
      20'h02678: out <= 12'h000;
      20'h02679: out <= 12'hc7f;
      20'h0267a: out <= 12'hfff;
      20'h0267b: out <= 12'hc7f;
      20'h0267c: out <= 12'h000;
      20'h0267d: out <= 12'h000;
      20'h0267e: out <= 12'h000;
      20'h0267f: out <= 12'h72f;
      20'h02680: out <= 12'hfff;
      20'h02681: out <= 12'h72f;
      20'h02682: out <= 12'h000;
      20'h02683: out <= 12'h000;
      20'h02684: out <= 12'h000;
      20'h02685: out <= 12'hc7f;
      20'h02686: out <= 12'hfff;
      20'h02687: out <= 12'hc7f;
      20'h02688: out <= 12'h222;
      20'h02689: out <= 12'h222;
      20'h0268a: out <= 12'h222;
      20'h0268b: out <= 12'h222;
      20'h0268c: out <= 12'h222;
      20'h0268d: out <= 12'h72f;
      20'h0268e: out <= 12'hfff;
      20'h0268f: out <= 12'hc7f;
      20'h02690: out <= 12'hc7f;
      20'h02691: out <= 12'hc7f;
      20'h02692: out <= 12'hc7f;
      20'h02693: out <= 12'hfff;
      20'h02694: out <= 12'h72f;
      20'h02695: out <= 12'h222;
      20'h02696: out <= 12'h222;
      20'h02697: out <= 12'h222;
      20'h02698: out <= 12'h000;
      20'h02699: out <= 12'h000;
      20'h0269a: out <= 12'h000;
      20'h0269b: out <= 12'h000;
      20'h0269c: out <= 12'h000;
      20'h0269d: out <= 12'h72f;
      20'h0269e: out <= 12'hfff;
      20'h0269f: out <= 12'hc7f;
      20'h026a0: out <= 12'hc7f;
      20'h026a1: out <= 12'hc7f;
      20'h026a2: out <= 12'hc7f;
      20'h026a3: out <= 12'hfff;
      20'h026a4: out <= 12'h72f;
      20'h026a5: out <= 12'h000;
      20'h026a6: out <= 12'h000;
      20'h026a7: out <= 12'h000;
      20'h026a8: out <= 12'h222;
      20'h026a9: out <= 12'hc7f;
      20'h026aa: out <= 12'hfff;
      20'h026ab: out <= 12'hc7f;
      20'h026ac: out <= 12'h72f;
      20'h026ad: out <= 12'hfff;
      20'h026ae: out <= 12'hc7f;
      20'h026af: out <= 12'hc7f;
      20'h026b0: out <= 12'hc7f;
      20'h026b1: out <= 12'hc7f;
      20'h026b2: out <= 12'hc7f;
      20'h026b3: out <= 12'hfff;
      20'h026b4: out <= 12'h72f;
      20'h026b5: out <= 12'hc7f;
      20'h026b6: out <= 12'hfff;
      20'h026b7: out <= 12'hc7f;
      20'h026b8: out <= 12'h000;
      20'h026b9: out <= 12'hc7f;
      20'h026ba: out <= 12'h72f;
      20'h026bb: out <= 12'hc7f;
      20'h026bc: out <= 12'h72f;
      20'h026bd: out <= 12'hfff;
      20'h026be: out <= 12'hc7f;
      20'h026bf: out <= 12'hc7f;
      20'h026c0: out <= 12'hc7f;
      20'h026c1: out <= 12'hc7f;
      20'h026c2: out <= 12'hc7f;
      20'h026c3: out <= 12'hfff;
      20'h026c4: out <= 12'h72f;
      20'h026c5: out <= 12'hc7f;
      20'h026c6: out <= 12'h72f;
      20'h026c7: out <= 12'hc7f;
      20'h026c8: out <= 12'h603;
      20'h026c9: out <= 12'h603;
      20'h026ca: out <= 12'h603;
      20'h026cb: out <= 12'h603;
      20'h026cc: out <= 12'h6af;
      20'h026cd: out <= 12'h4cd;
      20'h026ce: out <= 12'h4cd;
      20'h026cf: out <= 12'h6af;
      20'h026d0: out <= 12'hfff;
      20'h026d1: out <= 12'h4cd;
      20'h026d2: out <= 12'h4cd;
      20'h026d3: out <= 12'hfff;
      20'h026d4: out <= 12'h6af;
      20'h026d5: out <= 12'h4cd;
      20'h026d6: out <= 12'h4cd;
      20'h026d7: out <= 12'h6af;
      20'h026d8: out <= 12'hfff;
      20'h026d9: out <= 12'h4cd;
      20'h026da: out <= 12'h4cd;
      20'h026db: out <= 12'hfff;
      20'h026dc: out <= 12'h380;
      20'h026dd: out <= 12'hfff;
      20'h026de: out <= 12'h8d0;
      20'h026df: out <= 12'h8d0;
      20'h026e0: out <= 12'h380;
      20'h026e1: out <= 12'h000;
      20'h026e2: out <= 12'h8d0;
      20'h026e3: out <= 12'h000;
      20'h026e4: out <= 12'h380;
      20'h026e5: out <= 12'hfff;
      20'h026e6: out <= 12'h8d0;
      20'h026e7: out <= 12'h8d0;
      20'h026e8: out <= 12'h380;
      20'h026e9: out <= 12'h000;
      20'h026ea: out <= 12'h8d0;
      20'h026eb: out <= 12'h000;
      20'h026ec: out <= 12'h000;
      20'h026ed: out <= 12'h000;
      20'h026ee: out <= 12'hbbb;
      20'h026ef: out <= 12'hfff;
      20'h026f0: out <= 12'h000;
      20'h026f1: out <= 12'h000;
      20'h026f2: out <= 12'hbbb;
      20'h026f3: out <= 12'hfff;
      20'h026f4: out <= 12'h000;
      20'h026f5: out <= 12'h000;
      20'h026f6: out <= 12'hbbb;
      20'h026f7: out <= 12'hfff;
      20'h026f8: out <= 12'h000;
      20'h026f9: out <= 12'h000;
      20'h026fa: out <= 12'hbbb;
      20'h026fb: out <= 12'hfff;
      20'h026fc: out <= 12'h000;
      20'h026fd: out <= 12'h000;
      20'h026fe: out <= 12'h000;
      20'h026ff: out <= 12'h000;
      20'h02700: out <= 12'h000;
      20'h02701: out <= 12'h6af;
      20'h02702: out <= 12'h4cd;
      20'h02703: out <= 12'hfff;
      20'h02704: out <= 12'hfff;
      20'h02705: out <= 12'hfff;
      20'h02706: out <= 12'hfff;
      20'h02707: out <= 12'h4cd;
      20'h02708: out <= 12'h6af;
      20'h02709: out <= 12'h000;
      20'h0270a: out <= 12'h000;
      20'h0270b: out <= 12'h000;
      20'h0270c: out <= 12'h000;
      20'h0270d: out <= 12'h000;
      20'h0270e: out <= 12'h000;
      20'h0270f: out <= 12'h000;
      20'h02710: out <= 12'h000;
      20'h02711: out <= 12'h000;
      20'h02712: out <= 12'h000;
      20'h02713: out <= 12'h000;
      20'h02714: out <= 12'h000;
      20'h02715: out <= 12'h000;
      20'h02716: out <= 12'h000;
      20'h02717: out <= 12'h4cd;
      20'h02718: out <= 12'h4cd;
      20'h02719: out <= 12'hfff;
      20'h0271a: out <= 12'hfff;
      20'h0271b: out <= 12'h000;
      20'h0271c: out <= 12'h603;
      20'h0271d: out <= 12'h603;
      20'h0271e: out <= 12'h603;
      20'h0271f: out <= 12'h603;
      20'h02720: out <= 12'hee9;
      20'h02721: out <= 12'hf87;
      20'h02722: out <= 12'hee9;
      20'h02723: out <= 12'hf87;
      20'h02724: out <= 12'hf87;
      20'h02725: out <= 12'hb27;
      20'h02726: out <= 12'hf87;
      20'h02727: out <= 12'hb27;
      20'h02728: out <= 12'h000;
      20'h02729: out <= 12'h000;
      20'h0272a: out <= 12'h000;
      20'h0272b: out <= 12'h000;
      20'h0272c: out <= 12'h000;
      20'h0272d: out <= 12'h000;
      20'h0272e: out <= 12'h000;
      20'h0272f: out <= 12'h000;
      20'h02730: out <= 12'h000;
      20'h02731: out <= 12'h000;
      20'h02732: out <= 12'h000;
      20'h02733: out <= 12'h000;
      20'h02734: out <= 12'h000;
      20'h02735: out <= 12'h000;
      20'h02736: out <= 12'h000;
      20'h02737: out <= 12'h000;
      20'h02738: out <= 12'h916;
      20'h02739: out <= 12'h916;
      20'h0273a: out <= 12'h916;
      20'h0273b: out <= 12'h916;
      20'h0273c: out <= 12'h916;
      20'h0273d: out <= 12'h916;
      20'h0273e: out <= 12'h916;
      20'h0273f: out <= 12'h916;
      20'h02740: out <= 12'hd29;
      20'h02741: out <= 12'hd29;
      20'h02742: out <= 12'hd29;
      20'h02743: out <= 12'hd29;
      20'h02744: out <= 12'hd29;
      20'h02745: out <= 12'hd29;
      20'h02746: out <= 12'hd29;
      20'h02747: out <= 12'hd29;
      20'h02748: out <= 12'h000;
      20'h02749: out <= 12'h000;
      20'h0274a: out <= 12'h000;
      20'h0274b: out <= 12'h000;
      20'h0274c: out <= 12'h000;
      20'h0274d: out <= 12'h000;
      20'h0274e: out <= 12'h000;
      20'h0274f: out <= 12'h000;
      20'h02750: out <= 12'h000;
      20'h02751: out <= 12'h000;
      20'h02752: out <= 12'h000;
      20'h02753: out <= 12'h000;
      20'h02754: out <= 12'h000;
      20'h02755: out <= 12'h000;
      20'h02756: out <= 12'h000;
      20'h02757: out <= 12'h000;
      20'h02758: out <= 12'h000;
      20'h02759: out <= 12'h000;
      20'h0275a: out <= 12'h000;
      20'h0275b: out <= 12'h000;
      20'h0275c: out <= 12'h000;
      20'h0275d: out <= 12'h000;
      20'h0275e: out <= 12'h000;
      20'h0275f: out <= 12'h000;
      20'h02760: out <= 12'h222;
      20'h02761: out <= 12'h222;
      20'h02762: out <= 12'h72f;
      20'h02763: out <= 12'hfff;
      20'h02764: out <= 12'hc7f;
      20'h02765: out <= 12'hc7f;
      20'h02766: out <= 12'h72f;
      20'h02767: out <= 12'h72f;
      20'h02768: out <= 12'h72f;
      20'h02769: out <= 12'hc7f;
      20'h0276a: out <= 12'hfff;
      20'h0276b: out <= 12'h72f;
      20'h0276c: out <= 12'h222;
      20'h0276d: out <= 12'h222;
      20'h0276e: out <= 12'h222;
      20'h0276f: out <= 12'h222;
      20'h02770: out <= 12'h000;
      20'h02771: out <= 12'h000;
      20'h02772: out <= 12'h72f;
      20'h02773: out <= 12'hfff;
      20'h02774: out <= 12'hc7f;
      20'h02775: out <= 12'hc7f;
      20'h02776: out <= 12'h72f;
      20'h02777: out <= 12'h72f;
      20'h02778: out <= 12'h72f;
      20'h02779: out <= 12'hc7f;
      20'h0277a: out <= 12'hfff;
      20'h0277b: out <= 12'h72f;
      20'h0277c: out <= 12'h000;
      20'h0277d: out <= 12'h000;
      20'h0277e: out <= 12'h000;
      20'h0277f: out <= 12'h000;
      20'h02780: out <= 12'h222;
      20'h02781: out <= 12'hc7f;
      20'h02782: out <= 12'hfff;
      20'h02783: out <= 12'hc7f;
      20'h02784: out <= 12'h222;
      20'h02785: out <= 12'h72f;
      20'h02786: out <= 12'h72f;
      20'h02787: out <= 12'h72f;
      20'h02788: out <= 12'hfff;
      20'h02789: out <= 12'h72f;
      20'h0278a: out <= 12'h72f;
      20'h0278b: out <= 12'h72f;
      20'h0278c: out <= 12'h222;
      20'h0278d: out <= 12'hc7f;
      20'h0278e: out <= 12'hfff;
      20'h0278f: out <= 12'hc7f;
      20'h02790: out <= 12'h000;
      20'h02791: out <= 12'hc7f;
      20'h02792: out <= 12'h72f;
      20'h02793: out <= 12'hc7f;
      20'h02794: out <= 12'h000;
      20'h02795: out <= 12'h72f;
      20'h02796: out <= 12'h72f;
      20'h02797: out <= 12'h72f;
      20'h02798: out <= 12'hfff;
      20'h02799: out <= 12'h72f;
      20'h0279a: out <= 12'h72f;
      20'h0279b: out <= 12'h72f;
      20'h0279c: out <= 12'h000;
      20'h0279d: out <= 12'hc7f;
      20'h0279e: out <= 12'h72f;
      20'h0279f: out <= 12'hc7f;
      20'h027a0: out <= 12'h222;
      20'h027a1: out <= 12'h222;
      20'h027a2: out <= 12'h222;
      20'h027a3: out <= 12'h222;
      20'h027a4: out <= 12'h72f;
      20'h027a5: out <= 12'hfff;
      20'h027a6: out <= 12'hc7f;
      20'h027a7: out <= 12'h72f;
      20'h027a8: out <= 12'h72f;
      20'h027a9: out <= 12'h72f;
      20'h027aa: out <= 12'hc7f;
      20'h027ab: out <= 12'hc7f;
      20'h027ac: out <= 12'hfff;
      20'h027ad: out <= 12'h72f;
      20'h027ae: out <= 12'h222;
      20'h027af: out <= 12'h222;
      20'h027b0: out <= 12'h000;
      20'h027b1: out <= 12'h000;
      20'h027b2: out <= 12'h000;
      20'h027b3: out <= 12'h000;
      20'h027b4: out <= 12'h72f;
      20'h027b5: out <= 12'hfff;
      20'h027b6: out <= 12'hc7f;
      20'h027b7: out <= 12'h72f;
      20'h027b8: out <= 12'h72f;
      20'h027b9: out <= 12'h72f;
      20'h027ba: out <= 12'hc7f;
      20'h027bb: out <= 12'hc7f;
      20'h027bc: out <= 12'hfff;
      20'h027bd: out <= 12'h72f;
      20'h027be: out <= 12'h000;
      20'h027bf: out <= 12'h000;
      20'h027c0: out <= 12'h222;
      20'h027c1: out <= 12'hc7f;
      20'h027c2: out <= 12'h72f;
      20'h027c3: out <= 12'h72f;
      20'h027c4: out <= 12'hfff;
      20'h027c5: out <= 12'hc7f;
      20'h027c6: out <= 12'hc7f;
      20'h027c7: out <= 12'h72f;
      20'h027c8: out <= 12'h72f;
      20'h027c9: out <= 12'h72f;
      20'h027ca: out <= 12'hc7f;
      20'h027cb: out <= 12'hc7f;
      20'h027cc: out <= 12'hfff;
      20'h027cd: out <= 12'h72f;
      20'h027ce: out <= 12'h72f;
      20'h027cf: out <= 12'hc7f;
      20'h027d0: out <= 12'h000;
      20'h027d1: out <= 12'hc7f;
      20'h027d2: out <= 12'hfff;
      20'h027d3: out <= 12'h72f;
      20'h027d4: out <= 12'hfff;
      20'h027d5: out <= 12'hc7f;
      20'h027d6: out <= 12'hc7f;
      20'h027d7: out <= 12'h72f;
      20'h027d8: out <= 12'h72f;
      20'h027d9: out <= 12'h72f;
      20'h027da: out <= 12'hc7f;
      20'h027db: out <= 12'hc7f;
      20'h027dc: out <= 12'hfff;
      20'h027dd: out <= 12'h72f;
      20'h027de: out <= 12'hfff;
      20'h027df: out <= 12'hc7f;
      20'h027e0: out <= 12'h603;
      20'h027e1: out <= 12'h603;
      20'h027e2: out <= 12'h603;
      20'h027e3: out <= 12'h603;
      20'h027e4: out <= 12'hfff;
      20'h027e5: out <= 12'h6af;
      20'h027e6: out <= 12'h6af;
      20'h027e7: out <= 12'hfff;
      20'h027e8: out <= 12'h4cd;
      20'h027e9: out <= 12'h4cd;
      20'h027ea: out <= 12'h4cd;
      20'h027eb: out <= 12'h4cd;
      20'h027ec: out <= 12'hfff;
      20'h027ed: out <= 12'h6af;
      20'h027ee: out <= 12'h6af;
      20'h027ef: out <= 12'hfff;
      20'h027f0: out <= 12'h4cd;
      20'h027f1: out <= 12'h4cd;
      20'h027f2: out <= 12'h4cd;
      20'h027f3: out <= 12'h4cd;
      20'h027f4: out <= 12'hfff;
      20'h027f5: out <= 12'h8d0;
      20'h027f6: out <= 12'h8d0;
      20'h027f7: out <= 12'h380;
      20'h027f8: out <= 12'h8d0;
      20'h027f9: out <= 12'h8d0;
      20'h027fa: out <= 12'h000;
      20'h027fb: out <= 12'h380;
      20'h027fc: out <= 12'hfff;
      20'h027fd: out <= 12'h8d0;
      20'h027fe: out <= 12'h8d0;
      20'h027ff: out <= 12'h380;
      20'h02800: out <= 12'h8d0;
      20'h02801: out <= 12'h8d0;
      20'h02802: out <= 12'h000;
      20'h02803: out <= 12'h380;
      20'h02804: out <= 12'hfff;
      20'h02805: out <= 12'h666;
      20'h02806: out <= 12'h000;
      20'h02807: out <= 12'h000;
      20'h02808: out <= 12'hfff;
      20'h02809: out <= 12'h666;
      20'h0280a: out <= 12'h000;
      20'h0280b: out <= 12'h000;
      20'h0280c: out <= 12'hfff;
      20'h0280d: out <= 12'h666;
      20'h0280e: out <= 12'h000;
      20'h0280f: out <= 12'h000;
      20'h02810: out <= 12'hfff;
      20'h02811: out <= 12'h666;
      20'h02812: out <= 12'h000;
      20'h02813: out <= 12'h000;
      20'h02814: out <= 12'h000;
      20'h02815: out <= 12'h000;
      20'h02816: out <= 12'h000;
      20'h02817: out <= 12'h000;
      20'h02818: out <= 12'h000;
      20'h02819: out <= 12'h000;
      20'h0281a: out <= 12'h000;
      20'h0281b: out <= 12'h000;
      20'h0281c: out <= 12'h000;
      20'h0281d: out <= 12'h000;
      20'h0281e: out <= 12'h000;
      20'h0281f: out <= 12'h000;
      20'h02820: out <= 12'h000;
      20'h02821: out <= 12'h000;
      20'h02822: out <= 12'h000;
      20'h02823: out <= 12'h000;
      20'h02824: out <= 12'h000;
      20'h02825: out <= 12'h000;
      20'h02826: out <= 12'h000;
      20'h02827: out <= 12'h000;
      20'h02828: out <= 12'h000;
      20'h02829: out <= 12'h000;
      20'h0282a: out <= 12'h000;
      20'h0282b: out <= 12'h000;
      20'h0282c: out <= 12'h000;
      20'h0282d: out <= 12'h000;
      20'h0282e: out <= 12'h4cd;
      20'h0282f: out <= 12'h000;
      20'h02830: out <= 12'hfff;
      20'h02831: out <= 12'hfff;
      20'h02832: out <= 12'h4cd;
      20'h02833: out <= 12'h000;
      20'h02834: out <= 12'h603;
      20'h02835: out <= 12'h603;
      20'h02836: out <= 12'h603;
      20'h02837: out <= 12'h603;
      20'h02838: out <= 12'hee9;
      20'h02839: out <= 12'hf87;
      20'h0283a: out <= 12'hee9;
      20'h0283b: out <= 12'hf87;
      20'h0283c: out <= 12'hf87;
      20'h0283d: out <= 12'hb27;
      20'h0283e: out <= 12'hf87;
      20'h0283f: out <= 12'hb27;
      20'h02840: out <= 12'h000;
      20'h02841: out <= 12'h000;
      20'h02842: out <= 12'h000;
      20'h02843: out <= 12'h000;
      20'h02844: out <= 12'h000;
      20'h02845: out <= 12'h000;
      20'h02846: out <= 12'h000;
      20'h02847: out <= 12'h000;
      20'h02848: out <= 12'h000;
      20'h02849: out <= 12'h000;
      20'h0284a: out <= 12'h000;
      20'h0284b: out <= 12'h000;
      20'h0284c: out <= 12'h000;
      20'h0284d: out <= 12'h000;
      20'h0284e: out <= 12'h000;
      20'h0284f: out <= 12'h000;
      20'h02850: out <= 12'h916;
      20'h02851: out <= 12'h916;
      20'h02852: out <= 12'h916;
      20'h02853: out <= 12'h916;
      20'h02854: out <= 12'h916;
      20'h02855: out <= 12'h916;
      20'h02856: out <= 12'h916;
      20'h02857: out <= 12'h916;
      20'h02858: out <= 12'hd29;
      20'h02859: out <= 12'hd29;
      20'h0285a: out <= 12'hd29;
      20'h0285b: out <= 12'hd29;
      20'h0285c: out <= 12'hd29;
      20'h0285d: out <= 12'hd29;
      20'h0285e: out <= 12'hd29;
      20'h0285f: out <= 12'hd29;
      20'h02860: out <= 12'h000;
      20'h02861: out <= 12'h000;
      20'h02862: out <= 12'h000;
      20'h02863: out <= 12'h000;
      20'h02864: out <= 12'h000;
      20'h02865: out <= 12'h000;
      20'h02866: out <= 12'h000;
      20'h02867: out <= 12'h000;
      20'h02868: out <= 12'h000;
      20'h02869: out <= 12'h000;
      20'h0286a: out <= 12'h000;
      20'h0286b: out <= 12'h000;
      20'h0286c: out <= 12'h000;
      20'h0286d: out <= 12'h000;
      20'h0286e: out <= 12'h000;
      20'h0286f: out <= 12'h000;
      20'h02870: out <= 12'h000;
      20'h02871: out <= 12'h000;
      20'h02872: out <= 12'h000;
      20'h02873: out <= 12'h000;
      20'h02874: out <= 12'h000;
      20'h02875: out <= 12'h000;
      20'h02876: out <= 12'h000;
      20'h02877: out <= 12'h000;
      20'h02878: out <= 12'h222;
      20'h02879: out <= 12'h222;
      20'h0287a: out <= 12'h72f;
      20'h0287b: out <= 12'hc7f;
      20'h0287c: out <= 12'hc7f;
      20'h0287d: out <= 12'h72f;
      20'h0287e: out <= 12'h72f;
      20'h0287f: out <= 12'hc7f;
      20'h02880: out <= 12'h72f;
      20'h02881: out <= 12'h72f;
      20'h02882: out <= 12'hc7f;
      20'h02883: out <= 12'h72f;
      20'h02884: out <= 12'h222;
      20'h02885: out <= 12'h222;
      20'h02886: out <= 12'h222;
      20'h02887: out <= 12'h222;
      20'h02888: out <= 12'h000;
      20'h02889: out <= 12'h000;
      20'h0288a: out <= 12'h72f;
      20'h0288b: out <= 12'hc7f;
      20'h0288c: out <= 12'hc7f;
      20'h0288d: out <= 12'h72f;
      20'h0288e: out <= 12'h72f;
      20'h0288f: out <= 12'hc7f;
      20'h02890: out <= 12'h72f;
      20'h02891: out <= 12'h72f;
      20'h02892: out <= 12'hc7f;
      20'h02893: out <= 12'h72f;
      20'h02894: out <= 12'h000;
      20'h02895: out <= 12'h000;
      20'h02896: out <= 12'h000;
      20'h02897: out <= 12'h000;
      20'h02898: out <= 12'h222;
      20'h02899: out <= 12'hc7f;
      20'h0289a: out <= 12'h72f;
      20'h0289b: out <= 12'h72f;
      20'h0289c: out <= 12'h72f;
      20'h0289d: out <= 12'hfff;
      20'h0289e: out <= 12'hc7f;
      20'h0289f: out <= 12'h72f;
      20'h028a0: out <= 12'h72f;
      20'h028a1: out <= 12'h72f;
      20'h028a2: out <= 12'hc7f;
      20'h028a3: out <= 12'hfff;
      20'h028a4: out <= 12'h72f;
      20'h028a5: out <= 12'h72f;
      20'h028a6: out <= 12'h72f;
      20'h028a7: out <= 12'hc7f;
      20'h028a8: out <= 12'h000;
      20'h028a9: out <= 12'hc7f;
      20'h028aa: out <= 12'hfff;
      20'h028ab: out <= 12'h72f;
      20'h028ac: out <= 12'h72f;
      20'h028ad: out <= 12'hfff;
      20'h028ae: out <= 12'hc7f;
      20'h028af: out <= 12'h72f;
      20'h028b0: out <= 12'h72f;
      20'h028b1: out <= 12'h72f;
      20'h028b2: out <= 12'hc7f;
      20'h028b3: out <= 12'hfff;
      20'h028b4: out <= 12'h72f;
      20'h028b5: out <= 12'h72f;
      20'h028b6: out <= 12'hfff;
      20'h028b7: out <= 12'hc7f;
      20'h028b8: out <= 12'h222;
      20'h028b9: out <= 12'h222;
      20'h028ba: out <= 12'h222;
      20'h028bb: out <= 12'h222;
      20'h028bc: out <= 12'h72f;
      20'h028bd: out <= 12'hc7f;
      20'h028be: out <= 12'h72f;
      20'h028bf: out <= 12'h72f;
      20'h028c0: out <= 12'hc7f;
      20'h028c1: out <= 12'h72f;
      20'h028c2: out <= 12'h72f;
      20'h028c3: out <= 12'hc7f;
      20'h028c4: out <= 12'hc7f;
      20'h028c5: out <= 12'h72f;
      20'h028c6: out <= 12'h222;
      20'h028c7: out <= 12'h222;
      20'h028c8: out <= 12'h000;
      20'h028c9: out <= 12'h000;
      20'h028ca: out <= 12'h000;
      20'h028cb: out <= 12'h000;
      20'h028cc: out <= 12'h72f;
      20'h028cd: out <= 12'hc7f;
      20'h028ce: out <= 12'h72f;
      20'h028cf: out <= 12'h72f;
      20'h028d0: out <= 12'hc7f;
      20'h028d1: out <= 12'h72f;
      20'h028d2: out <= 12'h72f;
      20'h028d3: out <= 12'hc7f;
      20'h028d4: out <= 12'hc7f;
      20'h028d5: out <= 12'h72f;
      20'h028d6: out <= 12'h000;
      20'h028d7: out <= 12'h000;
      20'h028d8: out <= 12'h222;
      20'h028d9: out <= 12'hc7f;
      20'h028da: out <= 12'hfff;
      20'h028db: out <= 12'h72f;
      20'h028dc: out <= 12'hc7f;
      20'h028dd: out <= 12'hc7f;
      20'h028de: out <= 12'h72f;
      20'h028df: out <= 12'h72f;
      20'h028e0: out <= 12'hc7f;
      20'h028e1: out <= 12'h72f;
      20'h028e2: out <= 12'h72f;
      20'h028e3: out <= 12'hc7f;
      20'h028e4: out <= 12'hc7f;
      20'h028e5: out <= 12'h72f;
      20'h028e6: out <= 12'hfff;
      20'h028e7: out <= 12'hc7f;
      20'h028e8: out <= 12'h000;
      20'h028e9: out <= 12'hc7f;
      20'h028ea: out <= 12'h72f;
      20'h028eb: out <= 12'h72f;
      20'h028ec: out <= 12'hc7f;
      20'h028ed: out <= 12'hc7f;
      20'h028ee: out <= 12'h72f;
      20'h028ef: out <= 12'h72f;
      20'h028f0: out <= 12'hc7f;
      20'h028f1: out <= 12'h72f;
      20'h028f2: out <= 12'h72f;
      20'h028f3: out <= 12'hc7f;
      20'h028f4: out <= 12'hc7f;
      20'h028f5: out <= 12'h72f;
      20'h028f6: out <= 12'h72f;
      20'h028f7: out <= 12'hc7f;
      20'h028f8: out <= 12'h603;
      20'h028f9: out <= 12'h603;
      20'h028fa: out <= 12'h603;
      20'h028fb: out <= 12'h603;
      20'h028fc: out <= 12'h4cd;
      20'h028fd: out <= 12'hfff;
      20'h028fe: out <= 12'hfff;
      20'h028ff: out <= 12'h4cd;
      20'h02900: out <= 12'h4cd;
      20'h02901: out <= 12'h6af;
      20'h02902: out <= 12'h6af;
      20'h02903: out <= 12'h4cd;
      20'h02904: out <= 12'h4cd;
      20'h02905: out <= 12'hfff;
      20'h02906: out <= 12'hfff;
      20'h02907: out <= 12'h4cd;
      20'h02908: out <= 12'h4cd;
      20'h02909: out <= 12'h6af;
      20'h0290a: out <= 12'h6af;
      20'h0290b: out <= 12'h4cd;
      20'h0290c: out <= 12'h380;
      20'h0290d: out <= 12'h8d0;
      20'h0290e: out <= 12'h380;
      20'h0290f: out <= 12'h380;
      20'h02910: out <= 12'h8d0;
      20'h02911: out <= 12'h380;
      20'h02912: out <= 12'h380;
      20'h02913: out <= 12'h380;
      20'h02914: out <= 12'h380;
      20'h02915: out <= 12'h8d0;
      20'h02916: out <= 12'h380;
      20'h02917: out <= 12'h380;
      20'h02918: out <= 12'h8d0;
      20'h02919: out <= 12'h380;
      20'h0291a: out <= 12'h380;
      20'h0291b: out <= 12'h380;
      20'h0291c: out <= 12'hbbb;
      20'h0291d: out <= 12'hfff;
      20'h0291e: out <= 12'h000;
      20'h0291f: out <= 12'h000;
      20'h02920: out <= 12'hbbb;
      20'h02921: out <= 12'hfff;
      20'h02922: out <= 12'h000;
      20'h02923: out <= 12'h000;
      20'h02924: out <= 12'hbbb;
      20'h02925: out <= 12'hfff;
      20'h02926: out <= 12'h000;
      20'h02927: out <= 12'h000;
      20'h02928: out <= 12'hbbb;
      20'h02929: out <= 12'hfff;
      20'h0292a: out <= 12'h000;
      20'h0292b: out <= 12'h000;
      20'h0292c: out <= 12'h000;
      20'h0292d: out <= 12'h000;
      20'h0292e: out <= 12'h000;
      20'h0292f: out <= 12'h000;
      20'h02930: out <= 12'h6af;
      20'h02931: out <= 12'h000;
      20'h02932: out <= 12'h6af;
      20'h02933: out <= 12'h4cd;
      20'h02934: out <= 12'hfff;
      20'h02935: out <= 12'hfff;
      20'h02936: out <= 12'h4cd;
      20'h02937: out <= 12'h6af;
      20'h02938: out <= 12'h000;
      20'h02939: out <= 12'h000;
      20'h0293a: out <= 12'h000;
      20'h0293b: out <= 12'h000;
      20'h0293c: out <= 12'h000;
      20'h0293d: out <= 12'h000;
      20'h0293e: out <= 12'h000;
      20'h0293f: out <= 12'h000;
      20'h02940: out <= 12'h000;
      20'h02941: out <= 12'h000;
      20'h02942: out <= 12'h000;
      20'h02943: out <= 12'h000;
      20'h02944: out <= 12'h000;
      20'h02945: out <= 12'h4cd;
      20'h02946: out <= 12'h6af;
      20'h02947: out <= 12'hfff;
      20'h02948: out <= 12'h000;
      20'h02949: out <= 12'hfff;
      20'h0294a: out <= 12'h4cd;
      20'h0294b: out <= 12'h000;
      20'h0294c: out <= 12'h603;
      20'h0294d: out <= 12'h603;
      20'h0294e: out <= 12'h603;
      20'h0294f: out <= 12'h603;
      20'h02950: out <= 12'hee9;
      20'h02951: out <= 12'hf87;
      20'h02952: out <= 12'hee9;
      20'h02953: out <= 12'hb27;
      20'h02954: out <= 12'hb27;
      20'h02955: out <= 12'hb27;
      20'h02956: out <= 12'hf87;
      20'h02957: out <= 12'hb27;
      20'h02958: out <= 12'h000;
      20'h02959: out <= 12'h000;
      20'h0295a: out <= 12'h000;
      20'h0295b: out <= 12'h000;
      20'h0295c: out <= 12'h000;
      20'h0295d: out <= 12'h000;
      20'h0295e: out <= 12'h000;
      20'h0295f: out <= 12'h000;
      20'h02960: out <= 12'h000;
      20'h02961: out <= 12'h000;
      20'h02962: out <= 12'h000;
      20'h02963: out <= 12'h000;
      20'h02964: out <= 12'h000;
      20'h02965: out <= 12'h000;
      20'h02966: out <= 12'h000;
      20'h02967: out <= 12'h000;
      20'h02968: out <= 12'h916;
      20'h02969: out <= 12'h916;
      20'h0296a: out <= 12'h916;
      20'h0296b: out <= 12'h916;
      20'h0296c: out <= 12'h916;
      20'h0296d: out <= 12'h916;
      20'h0296e: out <= 12'h916;
      20'h0296f: out <= 12'h916;
      20'h02970: out <= 12'hd29;
      20'h02971: out <= 12'hd29;
      20'h02972: out <= 12'hd29;
      20'h02973: out <= 12'hd29;
      20'h02974: out <= 12'hd29;
      20'h02975: out <= 12'hd29;
      20'h02976: out <= 12'hd29;
      20'h02977: out <= 12'hd29;
      20'h02978: out <= 12'h000;
      20'h02979: out <= 12'h000;
      20'h0297a: out <= 12'h000;
      20'h0297b: out <= 12'h000;
      20'h0297c: out <= 12'h000;
      20'h0297d: out <= 12'h000;
      20'h0297e: out <= 12'h000;
      20'h0297f: out <= 12'h000;
      20'h02980: out <= 12'h000;
      20'h02981: out <= 12'h000;
      20'h02982: out <= 12'h000;
      20'h02983: out <= 12'h000;
      20'h02984: out <= 12'h000;
      20'h02985: out <= 12'h000;
      20'h02986: out <= 12'h000;
      20'h02987: out <= 12'h000;
      20'h02988: out <= 12'h000;
      20'h02989: out <= 12'h000;
      20'h0298a: out <= 12'h000;
      20'h0298b: out <= 12'h000;
      20'h0298c: out <= 12'h000;
      20'h0298d: out <= 12'h000;
      20'h0298e: out <= 12'h000;
      20'h0298f: out <= 12'h000;
      20'h02990: out <= 12'h222;
      20'h02991: out <= 12'h222;
      20'h02992: out <= 12'h72f;
      20'h02993: out <= 12'hc7f;
      20'h02994: out <= 12'h72f;
      20'h02995: out <= 12'h72f;
      20'h02996: out <= 12'hc7f;
      20'h02997: out <= 12'hfff;
      20'h02998: out <= 12'hc7f;
      20'h02999: out <= 12'h72f;
      20'h0299a: out <= 12'h72f;
      20'h0299b: out <= 12'h72f;
      20'h0299c: out <= 12'h72f;
      20'h0299d: out <= 12'h72f;
      20'h0299e: out <= 12'h72f;
      20'h0299f: out <= 12'hc7f;
      20'h029a0: out <= 12'h000;
      20'h029a1: out <= 12'h000;
      20'h029a2: out <= 12'h72f;
      20'h029a3: out <= 12'hc7f;
      20'h029a4: out <= 12'h72f;
      20'h029a5: out <= 12'h72f;
      20'h029a6: out <= 12'hc7f;
      20'h029a7: out <= 12'hfff;
      20'h029a8: out <= 12'hc7f;
      20'h029a9: out <= 12'h72f;
      20'h029aa: out <= 12'h72f;
      20'h029ab: out <= 12'h72f;
      20'h029ac: out <= 12'h72f;
      20'h029ad: out <= 12'h72f;
      20'h029ae: out <= 12'h72f;
      20'h029af: out <= 12'hc7f;
      20'h029b0: out <= 12'h222;
      20'h029b1: out <= 12'hc7f;
      20'h029b2: out <= 12'hfff;
      20'h029b3: out <= 12'h72f;
      20'h029b4: out <= 12'hfff;
      20'h029b5: out <= 12'hc7f;
      20'h029b6: out <= 12'h72f;
      20'h029b7: out <= 12'h72f;
      20'h029b8: out <= 12'hc7f;
      20'h029b9: out <= 12'h72f;
      20'h029ba: out <= 12'h72f;
      20'h029bb: out <= 12'hc7f;
      20'h029bc: out <= 12'hfff;
      20'h029bd: out <= 12'h72f;
      20'h029be: out <= 12'hfff;
      20'h029bf: out <= 12'hc7f;
      20'h029c0: out <= 12'h000;
      20'h029c1: out <= 12'hc7f;
      20'h029c2: out <= 12'h72f;
      20'h029c3: out <= 12'h72f;
      20'h029c4: out <= 12'hfff;
      20'h029c5: out <= 12'hc7f;
      20'h029c6: out <= 12'h72f;
      20'h029c7: out <= 12'h72f;
      20'h029c8: out <= 12'hc7f;
      20'h029c9: out <= 12'h72f;
      20'h029ca: out <= 12'h72f;
      20'h029cb: out <= 12'hc7f;
      20'h029cc: out <= 12'hfff;
      20'h029cd: out <= 12'h72f;
      20'h029ce: out <= 12'h72f;
      20'h029cf: out <= 12'hc7f;
      20'h029d0: out <= 12'hc7f;
      20'h029d1: out <= 12'h72f;
      20'h029d2: out <= 12'h72f;
      20'h029d3: out <= 12'h72f;
      20'h029d4: out <= 12'h72f;
      20'h029d5: out <= 12'h72f;
      20'h029d6: out <= 12'h72f;
      20'h029d7: out <= 12'hc7f;
      20'h029d8: out <= 12'hfff;
      20'h029d9: out <= 12'hc7f;
      20'h029da: out <= 12'h72f;
      20'h029db: out <= 12'h72f;
      20'h029dc: out <= 12'hc7f;
      20'h029dd: out <= 12'h72f;
      20'h029de: out <= 12'h222;
      20'h029df: out <= 12'h222;
      20'h029e0: out <= 12'hc7f;
      20'h029e1: out <= 12'h72f;
      20'h029e2: out <= 12'h72f;
      20'h029e3: out <= 12'h72f;
      20'h029e4: out <= 12'h72f;
      20'h029e5: out <= 12'h72f;
      20'h029e6: out <= 12'h72f;
      20'h029e7: out <= 12'hc7f;
      20'h029e8: out <= 12'hfff;
      20'h029e9: out <= 12'hc7f;
      20'h029ea: out <= 12'h72f;
      20'h029eb: out <= 12'h72f;
      20'h029ec: out <= 12'hc7f;
      20'h029ed: out <= 12'h72f;
      20'h029ee: out <= 12'h000;
      20'h029ef: out <= 12'h000;
      20'h029f0: out <= 12'h222;
      20'h029f1: out <= 12'hc7f;
      20'h029f2: out <= 12'h72f;
      20'h029f3: out <= 12'h72f;
      20'h029f4: out <= 12'hc7f;
      20'h029f5: out <= 12'h72f;
      20'h029f6: out <= 12'h72f;
      20'h029f7: out <= 12'hc7f;
      20'h029f8: out <= 12'hfff;
      20'h029f9: out <= 12'hc7f;
      20'h029fa: out <= 12'h72f;
      20'h029fb: out <= 12'h72f;
      20'h029fc: out <= 12'hc7f;
      20'h029fd: out <= 12'h72f;
      20'h029fe: out <= 12'h72f;
      20'h029ff: out <= 12'hc7f;
      20'h02a00: out <= 12'h000;
      20'h02a01: out <= 12'hc7f;
      20'h02a02: out <= 12'hfff;
      20'h02a03: out <= 12'h72f;
      20'h02a04: out <= 12'hc7f;
      20'h02a05: out <= 12'h72f;
      20'h02a06: out <= 12'h72f;
      20'h02a07: out <= 12'hc7f;
      20'h02a08: out <= 12'hfff;
      20'h02a09: out <= 12'hc7f;
      20'h02a0a: out <= 12'h72f;
      20'h02a0b: out <= 12'h72f;
      20'h02a0c: out <= 12'hc7f;
      20'h02a0d: out <= 12'h72f;
      20'h02a0e: out <= 12'hfff;
      20'h02a0f: out <= 12'hc7f;
      20'h02a10: out <= 12'h603;
      20'h02a11: out <= 12'h603;
      20'h02a12: out <= 12'h603;
      20'h02a13: out <= 12'h603;
      20'h02a14: out <= 12'h4cd;
      20'h02a15: out <= 12'h4cd;
      20'h02a16: out <= 12'h4cd;
      20'h02a17: out <= 12'h4cd;
      20'h02a18: out <= 12'h6af;
      20'h02a19: out <= 12'hfff;
      20'h02a1a: out <= 12'hfff;
      20'h02a1b: out <= 12'h6af;
      20'h02a1c: out <= 12'h4cd;
      20'h02a1d: out <= 12'h4cd;
      20'h02a1e: out <= 12'h4cd;
      20'h02a1f: out <= 12'h4cd;
      20'h02a20: out <= 12'h6af;
      20'h02a21: out <= 12'hfff;
      20'h02a22: out <= 12'hfff;
      20'h02a23: out <= 12'h6af;
      20'h02a24: out <= 12'h000;
      20'h02a25: out <= 12'h380;
      20'h02a26: out <= 12'h8d0;
      20'h02a27: out <= 12'h8d0;
      20'h02a28: out <= 12'h000;
      20'h02a29: out <= 12'h380;
      20'h02a2a: out <= 12'h000;
      20'h02a2b: out <= 12'h380;
      20'h02a2c: out <= 12'h000;
      20'h02a2d: out <= 12'h380;
      20'h02a2e: out <= 12'h8d0;
      20'h02a2f: out <= 12'h8d0;
      20'h02a30: out <= 12'h000;
      20'h02a31: out <= 12'h380;
      20'h02a32: out <= 12'h000;
      20'h02a33: out <= 12'h380;
      20'h02a34: out <= 12'h000;
      20'h02a35: out <= 12'h000;
      20'h02a36: out <= 12'hfff;
      20'h02a37: out <= 12'h666;
      20'h02a38: out <= 12'h000;
      20'h02a39: out <= 12'h000;
      20'h02a3a: out <= 12'hfff;
      20'h02a3b: out <= 12'h666;
      20'h02a3c: out <= 12'h000;
      20'h02a3d: out <= 12'h000;
      20'h02a3e: out <= 12'hfff;
      20'h02a3f: out <= 12'h666;
      20'h02a40: out <= 12'h000;
      20'h02a41: out <= 12'h000;
      20'h02a42: out <= 12'hfff;
      20'h02a43: out <= 12'h666;
      20'h02a44: out <= 12'h000;
      20'h02a45: out <= 12'h000;
      20'h02a46: out <= 12'h000;
      20'h02a47: out <= 12'h6af;
      20'h02a48: out <= 12'h4cd;
      20'h02a49: out <= 12'h000;
      20'h02a4a: out <= 12'h6af;
      20'h02a4b: out <= 12'h4cd;
      20'h02a4c: out <= 12'h000;
      20'h02a4d: out <= 12'h000;
      20'h02a4e: out <= 12'h4cd;
      20'h02a4f: out <= 12'h6af;
      20'h02a50: out <= 12'h000;
      20'h02a51: out <= 12'h000;
      20'h02a52: out <= 12'h000;
      20'h02a53: out <= 12'h000;
      20'h02a54: out <= 12'h000;
      20'h02a55: out <= 12'h000;
      20'h02a56: out <= 12'h6af;
      20'h02a57: out <= 12'h4cd;
      20'h02a58: out <= 12'h6af;
      20'h02a59: out <= 12'h000;
      20'h02a5a: out <= 12'h000;
      20'h02a5b: out <= 12'h000;
      20'h02a5c: out <= 12'h4cd;
      20'h02a5d: out <= 12'hfff;
      20'h02a5e: out <= 12'hfff;
      20'h02a5f: out <= 12'hfff;
      20'h02a60: out <= 12'h4cd;
      20'h02a61: out <= 12'h000;
      20'h02a62: out <= 12'h6af;
      20'h02a63: out <= 12'h000;
      20'h02a64: out <= 12'h603;
      20'h02a65: out <= 12'h603;
      20'h02a66: out <= 12'h603;
      20'h02a67: out <= 12'h603;
      20'h02a68: out <= 12'hee9;
      20'h02a69: out <= 12'hf87;
      20'h02a6a: out <= 12'hf87;
      20'h02a6b: out <= 12'hf87;
      20'h02a6c: out <= 12'hf87;
      20'h02a6d: out <= 12'hf87;
      20'h02a6e: out <= 12'hf87;
      20'h02a6f: out <= 12'hb27;
      20'h02a70: out <= 12'h000;
      20'h02a71: out <= 12'h000;
      20'h02a72: out <= 12'h000;
      20'h02a73: out <= 12'h000;
      20'h02a74: out <= 12'h000;
      20'h02a75: out <= 12'h000;
      20'h02a76: out <= 12'h000;
      20'h02a77: out <= 12'h000;
      20'h02a78: out <= 12'h000;
      20'h02a79: out <= 12'h000;
      20'h02a7a: out <= 12'h000;
      20'h02a7b: out <= 12'h000;
      20'h02a7c: out <= 12'h000;
      20'h02a7d: out <= 12'h000;
      20'h02a7e: out <= 12'h000;
      20'h02a7f: out <= 12'h000;
      20'h02a80: out <= 12'h916;
      20'h02a81: out <= 12'h916;
      20'h02a82: out <= 12'h916;
      20'h02a83: out <= 12'h916;
      20'h02a84: out <= 12'h916;
      20'h02a85: out <= 12'h916;
      20'h02a86: out <= 12'h916;
      20'h02a87: out <= 12'h916;
      20'h02a88: out <= 12'hd29;
      20'h02a89: out <= 12'hd29;
      20'h02a8a: out <= 12'hd29;
      20'h02a8b: out <= 12'hd29;
      20'h02a8c: out <= 12'hd29;
      20'h02a8d: out <= 12'hd29;
      20'h02a8e: out <= 12'hd29;
      20'h02a8f: out <= 12'hd29;
      20'h02a90: out <= 12'h000;
      20'h02a91: out <= 12'h000;
      20'h02a92: out <= 12'h000;
      20'h02a93: out <= 12'h000;
      20'h02a94: out <= 12'h000;
      20'h02a95: out <= 12'h000;
      20'h02a96: out <= 12'h000;
      20'h02a97: out <= 12'h000;
      20'h02a98: out <= 12'h000;
      20'h02a99: out <= 12'h000;
      20'h02a9a: out <= 12'h000;
      20'h02a9b: out <= 12'h000;
      20'h02a9c: out <= 12'h000;
      20'h02a9d: out <= 12'h000;
      20'h02a9e: out <= 12'h000;
      20'h02a9f: out <= 12'h000;
      20'h02aa0: out <= 12'h000;
      20'h02aa1: out <= 12'h000;
      20'h02aa2: out <= 12'h000;
      20'h02aa3: out <= 12'h000;
      20'h02aa4: out <= 12'h000;
      20'h02aa5: out <= 12'h000;
      20'h02aa6: out <= 12'h000;
      20'h02aa7: out <= 12'h000;
      20'h02aa8: out <= 12'h222;
      20'h02aa9: out <= 12'h222;
      20'h02aaa: out <= 12'h72f;
      20'h02aab: out <= 12'hc7f;
      20'h02aac: out <= 12'h72f;
      20'h02aad: out <= 12'hc7f;
      20'h02aae: out <= 12'hfff;
      20'h02aaf: out <= 12'hfff;
      20'h02ab0: out <= 12'hfff;
      20'h02ab1: out <= 12'hc7f;
      20'h02ab2: out <= 12'h72f;
      20'h02ab3: out <= 12'hfff;
      20'h02ab4: out <= 12'hfff;
      20'h02ab5: out <= 12'hfff;
      20'h02ab6: out <= 12'hfff;
      20'h02ab7: out <= 12'hfff;
      20'h02ab8: out <= 12'h000;
      20'h02ab9: out <= 12'h000;
      20'h02aba: out <= 12'h72f;
      20'h02abb: out <= 12'hc7f;
      20'h02abc: out <= 12'h72f;
      20'h02abd: out <= 12'hc7f;
      20'h02abe: out <= 12'hfff;
      20'h02abf: out <= 12'hfff;
      20'h02ac0: out <= 12'hfff;
      20'h02ac1: out <= 12'hc7f;
      20'h02ac2: out <= 12'h72f;
      20'h02ac3: out <= 12'hfff;
      20'h02ac4: out <= 12'hfff;
      20'h02ac5: out <= 12'hfff;
      20'h02ac6: out <= 12'hfff;
      20'h02ac7: out <= 12'hfff;
      20'h02ac8: out <= 12'h222;
      20'h02ac9: out <= 12'hc7f;
      20'h02aca: out <= 12'h72f;
      20'h02acb: out <= 12'h72f;
      20'h02acc: out <= 12'hc7f;
      20'h02acd: out <= 12'h72f;
      20'h02ace: out <= 12'h72f;
      20'h02acf: out <= 12'hc7f;
      20'h02ad0: out <= 12'hfff;
      20'h02ad1: out <= 12'hc7f;
      20'h02ad2: out <= 12'h72f;
      20'h02ad3: out <= 12'h72f;
      20'h02ad4: out <= 12'hc7f;
      20'h02ad5: out <= 12'h72f;
      20'h02ad6: out <= 12'h72f;
      20'h02ad7: out <= 12'hc7f;
      20'h02ad8: out <= 12'h000;
      20'h02ad9: out <= 12'hc7f;
      20'h02ada: out <= 12'hfff;
      20'h02adb: out <= 12'h72f;
      20'h02adc: out <= 12'hc7f;
      20'h02add: out <= 12'h72f;
      20'h02ade: out <= 12'h72f;
      20'h02adf: out <= 12'hc7f;
      20'h02ae0: out <= 12'hfff;
      20'h02ae1: out <= 12'hc7f;
      20'h02ae2: out <= 12'h72f;
      20'h02ae3: out <= 12'h72f;
      20'h02ae4: out <= 12'hc7f;
      20'h02ae5: out <= 12'h72f;
      20'h02ae6: out <= 12'hfff;
      20'h02ae7: out <= 12'hc7f;
      20'h02ae8: out <= 12'hfff;
      20'h02ae9: out <= 12'hfff;
      20'h02aea: out <= 12'hfff;
      20'h02aeb: out <= 12'hfff;
      20'h02aec: out <= 12'hfff;
      20'h02aed: out <= 12'h72f;
      20'h02aee: out <= 12'hc7f;
      20'h02aef: out <= 12'hfff;
      20'h02af0: out <= 12'hfff;
      20'h02af1: out <= 12'hfff;
      20'h02af2: out <= 12'hc7f;
      20'h02af3: out <= 12'h72f;
      20'h02af4: out <= 12'hc7f;
      20'h02af5: out <= 12'h72f;
      20'h02af6: out <= 12'h222;
      20'h02af7: out <= 12'h222;
      20'h02af8: out <= 12'hfff;
      20'h02af9: out <= 12'hfff;
      20'h02afa: out <= 12'hfff;
      20'h02afb: out <= 12'hfff;
      20'h02afc: out <= 12'hfff;
      20'h02afd: out <= 12'h72f;
      20'h02afe: out <= 12'hc7f;
      20'h02aff: out <= 12'hfff;
      20'h02b00: out <= 12'hfff;
      20'h02b01: out <= 12'hfff;
      20'h02b02: out <= 12'hc7f;
      20'h02b03: out <= 12'h72f;
      20'h02b04: out <= 12'hc7f;
      20'h02b05: out <= 12'h72f;
      20'h02b06: out <= 12'h000;
      20'h02b07: out <= 12'h000;
      20'h02b08: out <= 12'h222;
      20'h02b09: out <= 12'hc7f;
      20'h02b0a: out <= 12'hfff;
      20'h02b0b: out <= 12'h72f;
      20'h02b0c: out <= 12'hc7f;
      20'h02b0d: out <= 12'h72f;
      20'h02b0e: out <= 12'hc7f;
      20'h02b0f: out <= 12'hfff;
      20'h02b10: out <= 12'hfff;
      20'h02b11: out <= 12'hfff;
      20'h02b12: out <= 12'hc7f;
      20'h02b13: out <= 12'h72f;
      20'h02b14: out <= 12'hc7f;
      20'h02b15: out <= 12'h72f;
      20'h02b16: out <= 12'hfff;
      20'h02b17: out <= 12'hc7f;
      20'h02b18: out <= 12'h000;
      20'h02b19: out <= 12'hc7f;
      20'h02b1a: out <= 12'h72f;
      20'h02b1b: out <= 12'h72f;
      20'h02b1c: out <= 12'hc7f;
      20'h02b1d: out <= 12'h72f;
      20'h02b1e: out <= 12'hc7f;
      20'h02b1f: out <= 12'hfff;
      20'h02b20: out <= 12'hfff;
      20'h02b21: out <= 12'hfff;
      20'h02b22: out <= 12'hc7f;
      20'h02b23: out <= 12'h72f;
      20'h02b24: out <= 12'hc7f;
      20'h02b25: out <= 12'h72f;
      20'h02b26: out <= 12'h72f;
      20'h02b27: out <= 12'hc7f;
      20'h02b28: out <= 12'h603;
      20'h02b29: out <= 12'h603;
      20'h02b2a: out <= 12'h603;
      20'h02b2b: out <= 12'h603;
      20'h02b2c: out <= 12'h6af;
      20'h02b2d: out <= 12'h4cd;
      20'h02b2e: out <= 12'h4cd;
      20'h02b2f: out <= 12'h6af;
      20'h02b30: out <= 12'hfff;
      20'h02b31: out <= 12'h4cd;
      20'h02b32: out <= 12'h4cd;
      20'h02b33: out <= 12'hfff;
      20'h02b34: out <= 12'h6af;
      20'h02b35: out <= 12'h4cd;
      20'h02b36: out <= 12'h4cd;
      20'h02b37: out <= 12'h6af;
      20'h02b38: out <= 12'hfff;
      20'h02b39: out <= 12'h4cd;
      20'h02b3a: out <= 12'h4cd;
      20'h02b3b: out <= 12'hfff;
      20'h02b3c: out <= 12'h000;
      20'h02b3d: out <= 12'h000;
      20'h02b3e: out <= 12'h380;
      20'h02b3f: out <= 12'h380;
      20'h02b40: out <= 12'h380;
      20'h02b41: out <= 12'h380;
      20'h02b42: out <= 12'h000;
      20'h02b43: out <= 12'h000;
      20'h02b44: out <= 12'h000;
      20'h02b45: out <= 12'h000;
      20'h02b46: out <= 12'h380;
      20'h02b47: out <= 12'h380;
      20'h02b48: out <= 12'h380;
      20'h02b49: out <= 12'h380;
      20'h02b4a: out <= 12'h000;
      20'h02b4b: out <= 12'h000;
      20'h02b4c: out <= 12'h000;
      20'h02b4d: out <= 12'h000;
      20'h02b4e: out <= 12'hbbb;
      20'h02b4f: out <= 12'hfff;
      20'h02b50: out <= 12'h000;
      20'h02b51: out <= 12'h000;
      20'h02b52: out <= 12'hbbb;
      20'h02b53: out <= 12'hfff;
      20'h02b54: out <= 12'h000;
      20'h02b55: out <= 12'h000;
      20'h02b56: out <= 12'hbbb;
      20'h02b57: out <= 12'hfff;
      20'h02b58: out <= 12'h000;
      20'h02b59: out <= 12'h000;
      20'h02b5a: out <= 12'hbbb;
      20'h02b5b: out <= 12'hfff;
      20'h02b5c: out <= 12'h000;
      20'h02b5d: out <= 12'h000;
      20'h02b5e: out <= 12'h6af;
      20'h02b5f: out <= 12'h4cd;
      20'h02b60: out <= 12'hfff;
      20'h02b61: out <= 12'h000;
      20'h02b62: out <= 12'h6af;
      20'h02b63: out <= 12'h4cd;
      20'h02b64: out <= 12'h000;
      20'h02b65: out <= 12'h000;
      20'h02b66: out <= 12'h4cd;
      20'h02b67: out <= 12'h6af;
      20'h02b68: out <= 12'h000;
      20'h02b69: out <= 12'h000;
      20'h02b6a: out <= 12'h000;
      20'h02b6b: out <= 12'h000;
      20'h02b6c: out <= 12'h000;
      20'h02b6d: out <= 12'h000;
      20'h02b6e: out <= 12'h000;
      20'h02b6f: out <= 12'hfff;
      20'h02b70: out <= 12'hfff;
      20'h02b71: out <= 12'h000;
      20'h02b72: out <= 12'h000;
      20'h02b73: out <= 12'h6af;
      20'h02b74: out <= 12'hfff;
      20'h02b75: out <= 12'hfff;
      20'h02b76: out <= 12'hfff;
      20'h02b77: out <= 12'h4cd;
      20'h02b78: out <= 12'h6af;
      20'h02b79: out <= 12'h000;
      20'h02b7a: out <= 12'h000;
      20'h02b7b: out <= 12'h000;
      20'h02b7c: out <= 12'h603;
      20'h02b7d: out <= 12'h603;
      20'h02b7e: out <= 12'h603;
      20'h02b7f: out <= 12'h603;
      20'h02b80: out <= 12'hb27;
      20'h02b81: out <= 12'hb27;
      20'h02b82: out <= 12'hb27;
      20'h02b83: out <= 12'hb27;
      20'h02b84: out <= 12'hb27;
      20'h02b85: out <= 12'hb27;
      20'h02b86: out <= 12'hb27;
      20'h02b87: out <= 12'hb27;
      20'h02b88: out <= 12'h000;
      20'h02b89: out <= 12'h000;
      20'h02b8a: out <= 12'h000;
      20'h02b8b: out <= 12'h000;
      20'h02b8c: out <= 12'h000;
      20'h02b8d: out <= 12'h000;
      20'h02b8e: out <= 12'h000;
      20'h02b8f: out <= 12'h000;
      20'h02b90: out <= 12'h000;
      20'h02b91: out <= 12'h000;
      20'h02b92: out <= 12'h000;
      20'h02b93: out <= 12'h000;
      20'h02b94: out <= 12'h000;
      20'h02b95: out <= 12'h000;
      20'h02b96: out <= 12'h000;
      20'h02b97: out <= 12'h000;
      20'h02b98: out <= 12'h916;
      20'h02b99: out <= 12'h916;
      20'h02b9a: out <= 12'h916;
      20'h02b9b: out <= 12'h916;
      20'h02b9c: out <= 12'h916;
      20'h02b9d: out <= 12'h916;
      20'h02b9e: out <= 12'h916;
      20'h02b9f: out <= 12'h916;
      20'h02ba0: out <= 12'hd29;
      20'h02ba1: out <= 12'hd29;
      20'h02ba2: out <= 12'hd29;
      20'h02ba3: out <= 12'hd29;
      20'h02ba4: out <= 12'hd29;
      20'h02ba5: out <= 12'hd29;
      20'h02ba6: out <= 12'hd29;
      20'h02ba7: out <= 12'hd29;
      20'h02ba8: out <= 12'h000;
      20'h02ba9: out <= 12'h000;
      20'h02baa: out <= 12'h000;
      20'h02bab: out <= 12'h000;
      20'h02bac: out <= 12'h000;
      20'h02bad: out <= 12'h000;
      20'h02bae: out <= 12'h000;
      20'h02baf: out <= 12'h000;
      20'h02bb0: out <= 12'h000;
      20'h02bb1: out <= 12'h000;
      20'h02bb2: out <= 12'h000;
      20'h02bb3: out <= 12'h000;
      20'h02bb4: out <= 12'h000;
      20'h02bb5: out <= 12'h000;
      20'h02bb6: out <= 12'h000;
      20'h02bb7: out <= 12'h000;
      20'h02bb8: out <= 12'h000;
      20'h02bb9: out <= 12'h000;
      20'h02bba: out <= 12'h000;
      20'h02bbb: out <= 12'h000;
      20'h02bbc: out <= 12'h000;
      20'h02bbd: out <= 12'h000;
      20'h02bbe: out <= 12'h000;
      20'h02bbf: out <= 12'h000;
      20'h02bc0: out <= 12'h222;
      20'h02bc1: out <= 12'h222;
      20'h02bc2: out <= 12'h72f;
      20'h02bc3: out <= 12'hc7f;
      20'h02bc4: out <= 12'h72f;
      20'h02bc5: out <= 12'h72f;
      20'h02bc6: out <= 12'hc7f;
      20'h02bc7: out <= 12'hfff;
      20'h02bc8: out <= 12'hc7f;
      20'h02bc9: out <= 12'h72f;
      20'h02bca: out <= 12'h72f;
      20'h02bcb: out <= 12'h72f;
      20'h02bcc: out <= 12'h72f;
      20'h02bcd: out <= 12'h72f;
      20'h02bce: out <= 12'h72f;
      20'h02bcf: out <= 12'hc7f;
      20'h02bd0: out <= 12'h000;
      20'h02bd1: out <= 12'h000;
      20'h02bd2: out <= 12'h72f;
      20'h02bd3: out <= 12'hc7f;
      20'h02bd4: out <= 12'h72f;
      20'h02bd5: out <= 12'h72f;
      20'h02bd6: out <= 12'hc7f;
      20'h02bd7: out <= 12'hfff;
      20'h02bd8: out <= 12'hc7f;
      20'h02bd9: out <= 12'h72f;
      20'h02bda: out <= 12'h72f;
      20'h02bdb: out <= 12'h72f;
      20'h02bdc: out <= 12'h72f;
      20'h02bdd: out <= 12'h72f;
      20'h02bde: out <= 12'h72f;
      20'h02bdf: out <= 12'hc7f;
      20'h02be0: out <= 12'h222;
      20'h02be1: out <= 12'hc7f;
      20'h02be2: out <= 12'hfff;
      20'h02be3: out <= 12'h72f;
      20'h02be4: out <= 12'hc7f;
      20'h02be5: out <= 12'h72f;
      20'h02be6: out <= 12'hc7f;
      20'h02be7: out <= 12'hfff;
      20'h02be8: out <= 12'hfff;
      20'h02be9: out <= 12'hfff;
      20'h02bea: out <= 12'hc7f;
      20'h02beb: out <= 12'h72f;
      20'h02bec: out <= 12'hc7f;
      20'h02bed: out <= 12'h72f;
      20'h02bee: out <= 12'hfff;
      20'h02bef: out <= 12'hc7f;
      20'h02bf0: out <= 12'h000;
      20'h02bf1: out <= 12'hc7f;
      20'h02bf2: out <= 12'h72f;
      20'h02bf3: out <= 12'h72f;
      20'h02bf4: out <= 12'hc7f;
      20'h02bf5: out <= 12'h72f;
      20'h02bf6: out <= 12'hc7f;
      20'h02bf7: out <= 12'hfff;
      20'h02bf8: out <= 12'hfff;
      20'h02bf9: out <= 12'hfff;
      20'h02bfa: out <= 12'hc7f;
      20'h02bfb: out <= 12'h72f;
      20'h02bfc: out <= 12'hc7f;
      20'h02bfd: out <= 12'h72f;
      20'h02bfe: out <= 12'h72f;
      20'h02bff: out <= 12'hc7f;
      20'h02c00: out <= 12'hc7f;
      20'h02c01: out <= 12'h72f;
      20'h02c02: out <= 12'h72f;
      20'h02c03: out <= 12'h72f;
      20'h02c04: out <= 12'h72f;
      20'h02c05: out <= 12'h72f;
      20'h02c06: out <= 12'h72f;
      20'h02c07: out <= 12'hc7f;
      20'h02c08: out <= 12'hfff;
      20'h02c09: out <= 12'hc7f;
      20'h02c0a: out <= 12'h72f;
      20'h02c0b: out <= 12'h72f;
      20'h02c0c: out <= 12'hc7f;
      20'h02c0d: out <= 12'h72f;
      20'h02c0e: out <= 12'h222;
      20'h02c0f: out <= 12'h222;
      20'h02c10: out <= 12'hc7f;
      20'h02c11: out <= 12'h72f;
      20'h02c12: out <= 12'h72f;
      20'h02c13: out <= 12'h72f;
      20'h02c14: out <= 12'h72f;
      20'h02c15: out <= 12'h72f;
      20'h02c16: out <= 12'h72f;
      20'h02c17: out <= 12'hc7f;
      20'h02c18: out <= 12'hfff;
      20'h02c19: out <= 12'hc7f;
      20'h02c1a: out <= 12'h72f;
      20'h02c1b: out <= 12'h72f;
      20'h02c1c: out <= 12'hc7f;
      20'h02c1d: out <= 12'h72f;
      20'h02c1e: out <= 12'h000;
      20'h02c1f: out <= 12'h000;
      20'h02c20: out <= 12'h222;
      20'h02c21: out <= 12'hc7f;
      20'h02c22: out <= 12'h72f;
      20'h02c23: out <= 12'h72f;
      20'h02c24: out <= 12'hc7f;
      20'h02c25: out <= 12'h72f;
      20'h02c26: out <= 12'h72f;
      20'h02c27: out <= 12'hc7f;
      20'h02c28: out <= 12'hfff;
      20'h02c29: out <= 12'hc7f;
      20'h02c2a: out <= 12'h72f;
      20'h02c2b: out <= 12'h72f;
      20'h02c2c: out <= 12'hc7f;
      20'h02c2d: out <= 12'h72f;
      20'h02c2e: out <= 12'h72f;
      20'h02c2f: out <= 12'hc7f;
      20'h02c30: out <= 12'h000;
      20'h02c31: out <= 12'hc7f;
      20'h02c32: out <= 12'hfff;
      20'h02c33: out <= 12'h72f;
      20'h02c34: out <= 12'hc7f;
      20'h02c35: out <= 12'h72f;
      20'h02c36: out <= 12'h72f;
      20'h02c37: out <= 12'hc7f;
      20'h02c38: out <= 12'hfff;
      20'h02c39: out <= 12'hc7f;
      20'h02c3a: out <= 12'h72f;
      20'h02c3b: out <= 12'h72f;
      20'h02c3c: out <= 12'hc7f;
      20'h02c3d: out <= 12'h72f;
      20'h02c3e: out <= 12'hfff;
      20'h02c3f: out <= 12'hc7f;
      20'h02c40: out <= 12'h603;
      20'h02c41: out <= 12'h603;
      20'h02c42: out <= 12'h603;
      20'h02c43: out <= 12'h603;
      20'h02c44: out <= 12'hfff;
      20'h02c45: out <= 12'h6af;
      20'h02c46: out <= 12'h6af;
      20'h02c47: out <= 12'hfff;
      20'h02c48: out <= 12'h4cd;
      20'h02c49: out <= 12'h4cd;
      20'h02c4a: out <= 12'h4cd;
      20'h02c4b: out <= 12'h4cd;
      20'h02c4c: out <= 12'hfff;
      20'h02c4d: out <= 12'h6af;
      20'h02c4e: out <= 12'h6af;
      20'h02c4f: out <= 12'hfff;
      20'h02c50: out <= 12'h4cd;
      20'h02c51: out <= 12'h4cd;
      20'h02c52: out <= 12'h4cd;
      20'h02c53: out <= 12'h4cd;
      20'h02c54: out <= 12'h000;
      20'h02c55: out <= 12'h000;
      20'h02c56: out <= 12'hfff;
      20'h02c57: out <= 12'hfff;
      20'h02c58: out <= 12'hfff;
      20'h02c59: out <= 12'h8d0;
      20'h02c5a: out <= 12'h380;
      20'h02c5b: out <= 12'h000;
      20'h02c5c: out <= 12'h000;
      20'h02c5d: out <= 12'h000;
      20'h02c5e: out <= 12'hfff;
      20'h02c5f: out <= 12'hfff;
      20'h02c60: out <= 12'hfff;
      20'h02c61: out <= 12'h8d0;
      20'h02c62: out <= 12'h380;
      20'h02c63: out <= 12'h000;
      20'h02c64: out <= 12'hfff;
      20'h02c65: out <= 12'h666;
      20'h02c66: out <= 12'h000;
      20'h02c67: out <= 12'h000;
      20'h02c68: out <= 12'hfff;
      20'h02c69: out <= 12'h666;
      20'h02c6a: out <= 12'h000;
      20'h02c6b: out <= 12'h000;
      20'h02c6c: out <= 12'hfff;
      20'h02c6d: out <= 12'h666;
      20'h02c6e: out <= 12'h000;
      20'h02c6f: out <= 12'h000;
      20'h02c70: out <= 12'hfff;
      20'h02c71: out <= 12'h666;
      20'h02c72: out <= 12'h000;
      20'h02c73: out <= 12'h000;
      20'h02c74: out <= 12'h000;
      20'h02c75: out <= 12'h6af;
      20'h02c76: out <= 12'h4cd;
      20'h02c77: out <= 12'hfff;
      20'h02c78: out <= 12'hfff;
      20'h02c79: out <= 12'h000;
      20'h02c7a: out <= 12'h6af;
      20'h02c7b: out <= 12'h4cd;
      20'h02c7c: out <= 12'hfff;
      20'h02c7d: out <= 12'hfff;
      20'h02c7e: out <= 12'h4cd;
      20'h02c7f: out <= 12'h6af;
      20'h02c80: out <= 12'h000;
      20'h02c81: out <= 12'h000;
      20'h02c82: out <= 12'h000;
      20'h02c83: out <= 12'h000;
      20'h02c84: out <= 12'h000;
      20'h02c85: out <= 12'h000;
      20'h02c86: out <= 12'h6af;
      20'h02c87: out <= 12'h4cd;
      20'h02c88: out <= 12'h000;
      20'h02c89: out <= 12'h000;
      20'h02c8a: out <= 12'hfff;
      20'h02c8b: out <= 12'hfff;
      20'h02c8c: out <= 12'hfff;
      20'h02c8d: out <= 12'hfff;
      20'h02c8e: out <= 12'h4cd;
      20'h02c8f: out <= 12'h6af;
      20'h02c90: out <= 12'h000;
      20'h02c91: out <= 12'h000;
      20'h02c92: out <= 12'h4cd;
      20'h02c93: out <= 12'h000;
      20'h02c94: out <= 12'h603;
      20'h02c95: out <= 12'h603;
      20'h02c96: out <= 12'h603;
      20'h02c97: out <= 12'h603;
      20'h02c98: out <= 12'hee9;
      20'h02c99: out <= 12'hee9;
      20'h02c9a: out <= 12'hee9;
      20'h02c9b: out <= 12'hee9;
      20'h02c9c: out <= 12'hee9;
      20'h02c9d: out <= 12'hee9;
      20'h02c9e: out <= 12'hee9;
      20'h02c9f: out <= 12'hb27;
      20'h02ca0: out <= 12'h000;
      20'h02ca1: out <= 12'h000;
      20'h02ca2: out <= 12'h000;
      20'h02ca3: out <= 12'h000;
      20'h02ca4: out <= 12'h000;
      20'h02ca5: out <= 12'h000;
      20'h02ca6: out <= 12'h000;
      20'h02ca7: out <= 12'h000;
      20'h02ca8: out <= 12'h000;
      20'h02ca9: out <= 12'h000;
      20'h02caa: out <= 12'h000;
      20'h02cab: out <= 12'h000;
      20'h02cac: out <= 12'h000;
      20'h02cad: out <= 12'h000;
      20'h02cae: out <= 12'h000;
      20'h02caf: out <= 12'h000;
      20'h02cb0: out <= 12'h916;
      20'h02cb1: out <= 12'h916;
      20'h02cb2: out <= 12'h916;
      20'h02cb3: out <= 12'h916;
      20'h02cb4: out <= 12'h916;
      20'h02cb5: out <= 12'h916;
      20'h02cb6: out <= 12'h916;
      20'h02cb7: out <= 12'h916;
      20'h02cb8: out <= 12'hd29;
      20'h02cb9: out <= 12'hd29;
      20'h02cba: out <= 12'hd29;
      20'h02cbb: out <= 12'hd29;
      20'h02cbc: out <= 12'hd29;
      20'h02cbd: out <= 12'hd29;
      20'h02cbe: out <= 12'hd29;
      20'h02cbf: out <= 12'hd29;
      20'h02cc0: out <= 12'h000;
      20'h02cc1: out <= 12'h000;
      20'h02cc2: out <= 12'h000;
      20'h02cc3: out <= 12'h000;
      20'h02cc4: out <= 12'h000;
      20'h02cc5: out <= 12'h000;
      20'h02cc6: out <= 12'h000;
      20'h02cc7: out <= 12'h000;
      20'h02cc8: out <= 12'h000;
      20'h02cc9: out <= 12'h000;
      20'h02cca: out <= 12'h000;
      20'h02ccb: out <= 12'h000;
      20'h02ccc: out <= 12'h000;
      20'h02ccd: out <= 12'h000;
      20'h02cce: out <= 12'h000;
      20'h02ccf: out <= 12'h000;
      20'h02cd0: out <= 12'h000;
      20'h02cd1: out <= 12'h000;
      20'h02cd2: out <= 12'h000;
      20'h02cd3: out <= 12'h000;
      20'h02cd4: out <= 12'h000;
      20'h02cd5: out <= 12'h000;
      20'h02cd6: out <= 12'h000;
      20'h02cd7: out <= 12'h000;
      20'h02cd8: out <= 12'h222;
      20'h02cd9: out <= 12'h222;
      20'h02cda: out <= 12'h72f;
      20'h02cdb: out <= 12'hc7f;
      20'h02cdc: out <= 12'hc7f;
      20'h02cdd: out <= 12'h72f;
      20'h02cde: out <= 12'h72f;
      20'h02cdf: out <= 12'hc7f;
      20'h02ce0: out <= 12'h72f;
      20'h02ce1: out <= 12'h72f;
      20'h02ce2: out <= 12'hc7f;
      20'h02ce3: out <= 12'h72f;
      20'h02ce4: out <= 12'h222;
      20'h02ce5: out <= 12'h222;
      20'h02ce6: out <= 12'h222;
      20'h02ce7: out <= 12'h222;
      20'h02ce8: out <= 12'h000;
      20'h02ce9: out <= 12'h000;
      20'h02cea: out <= 12'h72f;
      20'h02ceb: out <= 12'hc7f;
      20'h02cec: out <= 12'hc7f;
      20'h02ced: out <= 12'h72f;
      20'h02cee: out <= 12'h72f;
      20'h02cef: out <= 12'hc7f;
      20'h02cf0: out <= 12'h72f;
      20'h02cf1: out <= 12'h72f;
      20'h02cf2: out <= 12'hc7f;
      20'h02cf3: out <= 12'h72f;
      20'h02cf4: out <= 12'h000;
      20'h02cf5: out <= 12'h000;
      20'h02cf6: out <= 12'h000;
      20'h02cf7: out <= 12'h000;
      20'h02cf8: out <= 12'h222;
      20'h02cf9: out <= 12'hc7f;
      20'h02cfa: out <= 12'h72f;
      20'h02cfb: out <= 12'h72f;
      20'h02cfc: out <= 12'hc7f;
      20'h02cfd: out <= 12'h72f;
      20'h02cfe: out <= 12'h72f;
      20'h02cff: out <= 12'hc7f;
      20'h02d00: out <= 12'hfff;
      20'h02d01: out <= 12'hc7f;
      20'h02d02: out <= 12'h72f;
      20'h02d03: out <= 12'h72f;
      20'h02d04: out <= 12'hc7f;
      20'h02d05: out <= 12'h72f;
      20'h02d06: out <= 12'h72f;
      20'h02d07: out <= 12'hc7f;
      20'h02d08: out <= 12'h000;
      20'h02d09: out <= 12'hc7f;
      20'h02d0a: out <= 12'hfff;
      20'h02d0b: out <= 12'h72f;
      20'h02d0c: out <= 12'hc7f;
      20'h02d0d: out <= 12'h72f;
      20'h02d0e: out <= 12'h72f;
      20'h02d0f: out <= 12'hc7f;
      20'h02d10: out <= 12'hfff;
      20'h02d11: out <= 12'hc7f;
      20'h02d12: out <= 12'h72f;
      20'h02d13: out <= 12'h72f;
      20'h02d14: out <= 12'hc7f;
      20'h02d15: out <= 12'h72f;
      20'h02d16: out <= 12'hfff;
      20'h02d17: out <= 12'hc7f;
      20'h02d18: out <= 12'h222;
      20'h02d19: out <= 12'h222;
      20'h02d1a: out <= 12'h222;
      20'h02d1b: out <= 12'h222;
      20'h02d1c: out <= 12'h72f;
      20'h02d1d: out <= 12'hc7f;
      20'h02d1e: out <= 12'h72f;
      20'h02d1f: out <= 12'h72f;
      20'h02d20: out <= 12'hc7f;
      20'h02d21: out <= 12'h72f;
      20'h02d22: out <= 12'h72f;
      20'h02d23: out <= 12'hc7f;
      20'h02d24: out <= 12'hc7f;
      20'h02d25: out <= 12'h72f;
      20'h02d26: out <= 12'h222;
      20'h02d27: out <= 12'h222;
      20'h02d28: out <= 12'h000;
      20'h02d29: out <= 12'h000;
      20'h02d2a: out <= 12'h000;
      20'h02d2b: out <= 12'h000;
      20'h02d2c: out <= 12'h72f;
      20'h02d2d: out <= 12'hc7f;
      20'h02d2e: out <= 12'h72f;
      20'h02d2f: out <= 12'h72f;
      20'h02d30: out <= 12'hc7f;
      20'h02d31: out <= 12'h72f;
      20'h02d32: out <= 12'h72f;
      20'h02d33: out <= 12'hc7f;
      20'h02d34: out <= 12'hc7f;
      20'h02d35: out <= 12'h72f;
      20'h02d36: out <= 12'h000;
      20'h02d37: out <= 12'h000;
      20'h02d38: out <= 12'h222;
      20'h02d39: out <= 12'hc7f;
      20'h02d3a: out <= 12'hfff;
      20'h02d3b: out <= 12'h72f;
      20'h02d3c: out <= 12'hfff;
      20'h02d3d: out <= 12'hc7f;
      20'h02d3e: out <= 12'h72f;
      20'h02d3f: out <= 12'h72f;
      20'h02d40: out <= 12'hc7f;
      20'h02d41: out <= 12'h72f;
      20'h02d42: out <= 12'h72f;
      20'h02d43: out <= 12'hc7f;
      20'h02d44: out <= 12'hfff;
      20'h02d45: out <= 12'h72f;
      20'h02d46: out <= 12'hfff;
      20'h02d47: out <= 12'hc7f;
      20'h02d48: out <= 12'h000;
      20'h02d49: out <= 12'hc7f;
      20'h02d4a: out <= 12'h72f;
      20'h02d4b: out <= 12'h72f;
      20'h02d4c: out <= 12'hfff;
      20'h02d4d: out <= 12'hc7f;
      20'h02d4e: out <= 12'h72f;
      20'h02d4f: out <= 12'h72f;
      20'h02d50: out <= 12'hc7f;
      20'h02d51: out <= 12'h72f;
      20'h02d52: out <= 12'h72f;
      20'h02d53: out <= 12'hc7f;
      20'h02d54: out <= 12'hfff;
      20'h02d55: out <= 12'h72f;
      20'h02d56: out <= 12'h72f;
      20'h02d57: out <= 12'hc7f;
      20'h02d58: out <= 12'h603;
      20'h02d59: out <= 12'h603;
      20'h02d5a: out <= 12'h603;
      20'h02d5b: out <= 12'h603;
      20'h02d5c: out <= 12'h4cd;
      20'h02d5d: out <= 12'hfff;
      20'h02d5e: out <= 12'hfff;
      20'h02d5f: out <= 12'h4cd;
      20'h02d60: out <= 12'h4cd;
      20'h02d61: out <= 12'h6af;
      20'h02d62: out <= 12'h6af;
      20'h02d63: out <= 12'h4cd;
      20'h02d64: out <= 12'h4cd;
      20'h02d65: out <= 12'hfff;
      20'h02d66: out <= 12'hfff;
      20'h02d67: out <= 12'h4cd;
      20'h02d68: out <= 12'h4cd;
      20'h02d69: out <= 12'h6af;
      20'h02d6a: out <= 12'h6af;
      20'h02d6b: out <= 12'h4cd;
      20'h02d6c: out <= 12'h000;
      20'h02d6d: out <= 12'hfff;
      20'h02d6e: out <= 12'h8d0;
      20'h02d6f: out <= 12'hfff;
      20'h02d70: out <= 12'h8d0;
      20'h02d71: out <= 12'h380;
      20'h02d72: out <= 12'h8d0;
      20'h02d73: out <= 12'h380;
      20'h02d74: out <= 12'h000;
      20'h02d75: out <= 12'hfff;
      20'h02d76: out <= 12'h8d0;
      20'h02d77: out <= 12'hfff;
      20'h02d78: out <= 12'h8d0;
      20'h02d79: out <= 12'h380;
      20'h02d7a: out <= 12'h8d0;
      20'h02d7b: out <= 12'h380;
      20'h02d7c: out <= 12'hbbb;
      20'h02d7d: out <= 12'hfff;
      20'h02d7e: out <= 12'h000;
      20'h02d7f: out <= 12'h000;
      20'h02d80: out <= 12'hbbb;
      20'h02d81: out <= 12'hfff;
      20'h02d82: out <= 12'h000;
      20'h02d83: out <= 12'h000;
      20'h02d84: out <= 12'hbbb;
      20'h02d85: out <= 12'hfff;
      20'h02d86: out <= 12'h000;
      20'h02d87: out <= 12'h000;
      20'h02d88: out <= 12'hbbb;
      20'h02d89: out <= 12'hfff;
      20'h02d8a: out <= 12'h000;
      20'h02d8b: out <= 12'h000;
      20'h02d8c: out <= 12'h000;
      20'h02d8d: out <= 12'h000;
      20'h02d8e: out <= 12'h000;
      20'h02d8f: out <= 12'h000;
      20'h02d90: out <= 12'h000;
      20'h02d91: out <= 12'h000;
      20'h02d92: out <= 12'h6af;
      20'h02d93: out <= 12'h4cd;
      20'h02d94: out <= 12'hfff;
      20'h02d95: out <= 12'h000;
      20'h02d96: out <= 12'h000;
      20'h02d97: out <= 12'h000;
      20'h02d98: out <= 12'h000;
      20'h02d99: out <= 12'h000;
      20'h02d9a: out <= 12'h000;
      20'h02d9b: out <= 12'h000;
      20'h02d9c: out <= 12'h000;
      20'h02d9d: out <= 12'h000;
      20'h02d9e: out <= 12'h6af;
      20'h02d9f: out <= 12'h000;
      20'h02da0: out <= 12'h000;
      20'h02da1: out <= 12'h4cd;
      20'h02da2: out <= 12'hfff;
      20'h02da3: out <= 12'hfff;
      20'h02da4: out <= 12'hfff;
      20'h02da5: out <= 12'h000;
      20'h02da6: out <= 12'h000;
      20'h02da7: out <= 12'h000;
      20'h02da8: out <= 12'h000;
      20'h02da9: out <= 12'h000;
      20'h02daa: out <= 12'h000;
      20'h02dab: out <= 12'h000;
      20'h02dac: out <= 12'h603;
      20'h02dad: out <= 12'h603;
      20'h02dae: out <= 12'h603;
      20'h02daf: out <= 12'h603;
      20'h02db0: out <= 12'hee9;
      20'h02db1: out <= 12'hf87;
      20'h02db2: out <= 12'hf87;
      20'h02db3: out <= 12'hf87;
      20'h02db4: out <= 12'hf87;
      20'h02db5: out <= 12'hf87;
      20'h02db6: out <= 12'hf87;
      20'h02db7: out <= 12'hb27;
      20'h02db8: out <= 12'h000;
      20'h02db9: out <= 12'h000;
      20'h02dba: out <= 12'h000;
      20'h02dbb: out <= 12'h000;
      20'h02dbc: out <= 12'h000;
      20'h02dbd: out <= 12'h000;
      20'h02dbe: out <= 12'h000;
      20'h02dbf: out <= 12'h000;
      20'h02dc0: out <= 12'h000;
      20'h02dc1: out <= 12'h000;
      20'h02dc2: out <= 12'h000;
      20'h02dc3: out <= 12'h000;
      20'h02dc4: out <= 12'h000;
      20'h02dc5: out <= 12'h000;
      20'h02dc6: out <= 12'h000;
      20'h02dc7: out <= 12'h000;
      20'h02dc8: out <= 12'h916;
      20'h02dc9: out <= 12'h916;
      20'h02dca: out <= 12'h916;
      20'h02dcb: out <= 12'h916;
      20'h02dcc: out <= 12'h916;
      20'h02dcd: out <= 12'h916;
      20'h02dce: out <= 12'h916;
      20'h02dcf: out <= 12'h916;
      20'h02dd0: out <= 12'hd29;
      20'h02dd1: out <= 12'hd29;
      20'h02dd2: out <= 12'hd29;
      20'h02dd3: out <= 12'hd29;
      20'h02dd4: out <= 12'hd29;
      20'h02dd5: out <= 12'hd29;
      20'h02dd6: out <= 12'hd29;
      20'h02dd7: out <= 12'hd29;
      20'h02dd8: out <= 12'h000;
      20'h02dd9: out <= 12'h000;
      20'h02dda: out <= 12'h000;
      20'h02ddb: out <= 12'h000;
      20'h02ddc: out <= 12'h000;
      20'h02ddd: out <= 12'h000;
      20'h02dde: out <= 12'h000;
      20'h02ddf: out <= 12'h000;
      20'h02de0: out <= 12'h000;
      20'h02de1: out <= 12'h000;
      20'h02de2: out <= 12'h000;
      20'h02de3: out <= 12'h000;
      20'h02de4: out <= 12'h000;
      20'h02de5: out <= 12'h000;
      20'h02de6: out <= 12'h000;
      20'h02de7: out <= 12'h000;
      20'h02de8: out <= 12'h000;
      20'h02de9: out <= 12'h000;
      20'h02dea: out <= 12'h000;
      20'h02deb: out <= 12'h000;
      20'h02dec: out <= 12'h000;
      20'h02ded: out <= 12'h000;
      20'h02dee: out <= 12'h000;
      20'h02def: out <= 12'h000;
      20'h02df0: out <= 12'h222;
      20'h02df1: out <= 12'h222;
      20'h02df2: out <= 12'h72f;
      20'h02df3: out <= 12'hfff;
      20'h02df4: out <= 12'hc7f;
      20'h02df5: out <= 12'hc7f;
      20'h02df6: out <= 12'h72f;
      20'h02df7: out <= 12'h72f;
      20'h02df8: out <= 12'h72f;
      20'h02df9: out <= 12'hc7f;
      20'h02dfa: out <= 12'hfff;
      20'h02dfb: out <= 12'h72f;
      20'h02dfc: out <= 12'h222;
      20'h02dfd: out <= 12'h222;
      20'h02dfe: out <= 12'h222;
      20'h02dff: out <= 12'h222;
      20'h02e00: out <= 12'h000;
      20'h02e01: out <= 12'h000;
      20'h02e02: out <= 12'h72f;
      20'h02e03: out <= 12'hfff;
      20'h02e04: out <= 12'hc7f;
      20'h02e05: out <= 12'hc7f;
      20'h02e06: out <= 12'h72f;
      20'h02e07: out <= 12'h72f;
      20'h02e08: out <= 12'h72f;
      20'h02e09: out <= 12'hc7f;
      20'h02e0a: out <= 12'hfff;
      20'h02e0b: out <= 12'h72f;
      20'h02e0c: out <= 12'h000;
      20'h02e0d: out <= 12'h000;
      20'h02e0e: out <= 12'h000;
      20'h02e0f: out <= 12'h000;
      20'h02e10: out <= 12'h222;
      20'h02e11: out <= 12'hc7f;
      20'h02e12: out <= 12'hfff;
      20'h02e13: out <= 12'h72f;
      20'h02e14: out <= 12'hc7f;
      20'h02e15: out <= 12'hc7f;
      20'h02e16: out <= 12'h72f;
      20'h02e17: out <= 12'h72f;
      20'h02e18: out <= 12'hc7f;
      20'h02e19: out <= 12'h72f;
      20'h02e1a: out <= 12'h72f;
      20'h02e1b: out <= 12'hc7f;
      20'h02e1c: out <= 12'hc7f;
      20'h02e1d: out <= 12'h72f;
      20'h02e1e: out <= 12'hfff;
      20'h02e1f: out <= 12'hc7f;
      20'h02e20: out <= 12'h000;
      20'h02e21: out <= 12'hc7f;
      20'h02e22: out <= 12'h72f;
      20'h02e23: out <= 12'h72f;
      20'h02e24: out <= 12'hc7f;
      20'h02e25: out <= 12'hc7f;
      20'h02e26: out <= 12'h72f;
      20'h02e27: out <= 12'h72f;
      20'h02e28: out <= 12'hc7f;
      20'h02e29: out <= 12'h72f;
      20'h02e2a: out <= 12'h72f;
      20'h02e2b: out <= 12'hc7f;
      20'h02e2c: out <= 12'hc7f;
      20'h02e2d: out <= 12'h72f;
      20'h02e2e: out <= 12'h72f;
      20'h02e2f: out <= 12'hc7f;
      20'h02e30: out <= 12'h222;
      20'h02e31: out <= 12'h222;
      20'h02e32: out <= 12'h222;
      20'h02e33: out <= 12'h222;
      20'h02e34: out <= 12'h72f;
      20'h02e35: out <= 12'hfff;
      20'h02e36: out <= 12'hc7f;
      20'h02e37: out <= 12'h72f;
      20'h02e38: out <= 12'h72f;
      20'h02e39: out <= 12'h72f;
      20'h02e3a: out <= 12'hc7f;
      20'h02e3b: out <= 12'hc7f;
      20'h02e3c: out <= 12'hfff;
      20'h02e3d: out <= 12'h72f;
      20'h02e3e: out <= 12'h222;
      20'h02e3f: out <= 12'h222;
      20'h02e40: out <= 12'h000;
      20'h02e41: out <= 12'h000;
      20'h02e42: out <= 12'h000;
      20'h02e43: out <= 12'h000;
      20'h02e44: out <= 12'h72f;
      20'h02e45: out <= 12'hfff;
      20'h02e46: out <= 12'hc7f;
      20'h02e47: out <= 12'h72f;
      20'h02e48: out <= 12'h72f;
      20'h02e49: out <= 12'h72f;
      20'h02e4a: out <= 12'hc7f;
      20'h02e4b: out <= 12'hc7f;
      20'h02e4c: out <= 12'hfff;
      20'h02e4d: out <= 12'h72f;
      20'h02e4e: out <= 12'h000;
      20'h02e4f: out <= 12'h000;
      20'h02e50: out <= 12'h222;
      20'h02e51: out <= 12'hc7f;
      20'h02e52: out <= 12'h72f;
      20'h02e53: out <= 12'h72f;
      20'h02e54: out <= 12'h72f;
      20'h02e55: out <= 12'hfff;
      20'h02e56: out <= 12'hc7f;
      20'h02e57: out <= 12'h72f;
      20'h02e58: out <= 12'h72f;
      20'h02e59: out <= 12'h72f;
      20'h02e5a: out <= 12'hc7f;
      20'h02e5b: out <= 12'hfff;
      20'h02e5c: out <= 12'h72f;
      20'h02e5d: out <= 12'h72f;
      20'h02e5e: out <= 12'h72f;
      20'h02e5f: out <= 12'hc7f;
      20'h02e60: out <= 12'h000;
      20'h02e61: out <= 12'hc7f;
      20'h02e62: out <= 12'hfff;
      20'h02e63: out <= 12'h72f;
      20'h02e64: out <= 12'h72f;
      20'h02e65: out <= 12'hfff;
      20'h02e66: out <= 12'hc7f;
      20'h02e67: out <= 12'h72f;
      20'h02e68: out <= 12'h72f;
      20'h02e69: out <= 12'h72f;
      20'h02e6a: out <= 12'hc7f;
      20'h02e6b: out <= 12'hfff;
      20'h02e6c: out <= 12'h72f;
      20'h02e6d: out <= 12'h72f;
      20'h02e6e: out <= 12'hfff;
      20'h02e6f: out <= 12'hc7f;
      20'h02e70: out <= 12'h603;
      20'h02e71: out <= 12'h603;
      20'h02e72: out <= 12'h603;
      20'h02e73: out <= 12'h603;
      20'h02e74: out <= 12'h4cd;
      20'h02e75: out <= 12'h4cd;
      20'h02e76: out <= 12'h4cd;
      20'h02e77: out <= 12'h4cd;
      20'h02e78: out <= 12'h6af;
      20'h02e79: out <= 12'hfff;
      20'h02e7a: out <= 12'hfff;
      20'h02e7b: out <= 12'h6af;
      20'h02e7c: out <= 12'h4cd;
      20'h02e7d: out <= 12'h4cd;
      20'h02e7e: out <= 12'h4cd;
      20'h02e7f: out <= 12'h4cd;
      20'h02e80: out <= 12'h6af;
      20'h02e81: out <= 12'hfff;
      20'h02e82: out <= 12'hfff;
      20'h02e83: out <= 12'h6af;
      20'h02e84: out <= 12'hfff;
      20'h02e85: out <= 12'h8d0;
      20'h02e86: out <= 12'hfff;
      20'h02e87: out <= 12'h8d0;
      20'h02e88: out <= 12'h8d0;
      20'h02e89: out <= 12'h8d0;
      20'h02e8a: out <= 12'h380;
      20'h02e8b: out <= 12'h8d0;
      20'h02e8c: out <= 12'hfff;
      20'h02e8d: out <= 12'h8d0;
      20'h02e8e: out <= 12'hfff;
      20'h02e8f: out <= 12'h8d0;
      20'h02e90: out <= 12'h8d0;
      20'h02e91: out <= 12'h8d0;
      20'h02e92: out <= 12'h380;
      20'h02e93: out <= 12'h8d0;
      20'h02e94: out <= 12'h000;
      20'h02e95: out <= 12'h000;
      20'h02e96: out <= 12'hfff;
      20'h02e97: out <= 12'h666;
      20'h02e98: out <= 12'h000;
      20'h02e99: out <= 12'h000;
      20'h02e9a: out <= 12'hfff;
      20'h02e9b: out <= 12'h666;
      20'h02e9c: out <= 12'h000;
      20'h02e9d: out <= 12'h000;
      20'h02e9e: out <= 12'hfff;
      20'h02e9f: out <= 12'h666;
      20'h02ea0: out <= 12'h000;
      20'h02ea1: out <= 12'h000;
      20'h02ea2: out <= 12'hfff;
      20'h02ea3: out <= 12'h666;
      20'h02ea4: out <= 12'h000;
      20'h02ea5: out <= 12'h6af;
      20'h02ea6: out <= 12'h4cd;
      20'h02ea7: out <= 12'hfff;
      20'h02ea8: out <= 12'hfff;
      20'h02ea9: out <= 12'h000;
      20'h02eaa: out <= 12'h6af;
      20'h02eab: out <= 12'h4cd;
      20'h02eac: out <= 12'hfff;
      20'h02ead: out <= 12'h000;
      20'h02eae: out <= 12'h6af;
      20'h02eaf: out <= 12'h4cd;
      20'h02eb0: out <= 12'hfff;
      20'h02eb1: out <= 12'hfff;
      20'h02eb2: out <= 12'h4cd;
      20'h02eb3: out <= 12'h6af;
      20'h02eb4: out <= 12'h000;
      20'h02eb5: out <= 12'h000;
      20'h02eb6: out <= 12'h000;
      20'h02eb7: out <= 12'hfff;
      20'h02eb8: out <= 12'h000;
      20'h02eb9: out <= 12'h000;
      20'h02eba: out <= 12'hfff;
      20'h02ebb: out <= 12'h4cd;
      20'h02ebc: out <= 12'h000;
      20'h02ebd: out <= 12'h6af;
      20'h02ebe: out <= 12'h4cd;
      20'h02ebf: out <= 12'h4cd;
      20'h02ec0: out <= 12'h4cd;
      20'h02ec1: out <= 12'h6af;
      20'h02ec2: out <= 12'h000;
      20'h02ec3: out <= 12'h000;
      20'h02ec4: out <= 12'h603;
      20'h02ec5: out <= 12'h603;
      20'h02ec6: out <= 12'h603;
      20'h02ec7: out <= 12'h603;
      20'h02ec8: out <= 12'hee9;
      20'h02ec9: out <= 12'hf87;
      20'h02eca: out <= 12'hee9;
      20'h02ecb: out <= 12'hee9;
      20'h02ecc: out <= 12'hee9;
      20'h02ecd: out <= 12'hb27;
      20'h02ece: out <= 12'hf87;
      20'h02ecf: out <= 12'hb27;
      20'h02ed0: out <= 12'h000;
      20'h02ed1: out <= 12'h000;
      20'h02ed2: out <= 12'h000;
      20'h02ed3: out <= 12'h000;
      20'h02ed4: out <= 12'h000;
      20'h02ed5: out <= 12'h000;
      20'h02ed6: out <= 12'h000;
      20'h02ed7: out <= 12'h000;
      20'h02ed8: out <= 12'h000;
      20'h02ed9: out <= 12'h000;
      20'h02eda: out <= 12'h000;
      20'h02edb: out <= 12'h000;
      20'h02edc: out <= 12'h000;
      20'h02edd: out <= 12'h000;
      20'h02ede: out <= 12'h000;
      20'h02edf: out <= 12'h000;
      20'h02ee0: out <= 12'h916;
      20'h02ee1: out <= 12'h916;
      20'h02ee2: out <= 12'h916;
      20'h02ee3: out <= 12'h916;
      20'h02ee4: out <= 12'h916;
      20'h02ee5: out <= 12'h916;
      20'h02ee6: out <= 12'h916;
      20'h02ee7: out <= 12'h916;
      20'h02ee8: out <= 12'hd29;
      20'h02ee9: out <= 12'hd29;
      20'h02eea: out <= 12'hd29;
      20'h02eeb: out <= 12'hd29;
      20'h02eec: out <= 12'hd29;
      20'h02eed: out <= 12'hd29;
      20'h02eee: out <= 12'hd29;
      20'h02eef: out <= 12'hd29;
      20'h02ef0: out <= 12'h000;
      20'h02ef1: out <= 12'h000;
      20'h02ef2: out <= 12'h000;
      20'h02ef3: out <= 12'h000;
      20'h02ef4: out <= 12'h000;
      20'h02ef5: out <= 12'h000;
      20'h02ef6: out <= 12'h000;
      20'h02ef7: out <= 12'h000;
      20'h02ef8: out <= 12'h000;
      20'h02ef9: out <= 12'h000;
      20'h02efa: out <= 12'h000;
      20'h02efb: out <= 12'h000;
      20'h02efc: out <= 12'h000;
      20'h02efd: out <= 12'h000;
      20'h02efe: out <= 12'h000;
      20'h02eff: out <= 12'h000;
      20'h02f00: out <= 12'h000;
      20'h02f01: out <= 12'h000;
      20'h02f02: out <= 12'h000;
      20'h02f03: out <= 12'h000;
      20'h02f04: out <= 12'h000;
      20'h02f05: out <= 12'h000;
      20'h02f06: out <= 12'h000;
      20'h02f07: out <= 12'h000;
      20'h02f08: out <= 12'h222;
      20'h02f09: out <= 12'h222;
      20'h02f0a: out <= 12'h222;
      20'h02f0b: out <= 12'h72f;
      20'h02f0c: out <= 12'hfff;
      20'h02f0d: out <= 12'hc7f;
      20'h02f0e: out <= 12'hc7f;
      20'h02f0f: out <= 12'hc7f;
      20'h02f10: out <= 12'hc7f;
      20'h02f11: out <= 12'hfff;
      20'h02f12: out <= 12'h72f;
      20'h02f13: out <= 12'h222;
      20'h02f14: out <= 12'h222;
      20'h02f15: out <= 12'h222;
      20'h02f16: out <= 12'h222;
      20'h02f17: out <= 12'h222;
      20'h02f18: out <= 12'h000;
      20'h02f19: out <= 12'h000;
      20'h02f1a: out <= 12'h000;
      20'h02f1b: out <= 12'h72f;
      20'h02f1c: out <= 12'hfff;
      20'h02f1d: out <= 12'hc7f;
      20'h02f1e: out <= 12'hc7f;
      20'h02f1f: out <= 12'hc7f;
      20'h02f20: out <= 12'hc7f;
      20'h02f21: out <= 12'hfff;
      20'h02f22: out <= 12'h72f;
      20'h02f23: out <= 12'h000;
      20'h02f24: out <= 12'h000;
      20'h02f25: out <= 12'h000;
      20'h02f26: out <= 12'h000;
      20'h02f27: out <= 12'h000;
      20'h02f28: out <= 12'h222;
      20'h02f29: out <= 12'hc7f;
      20'h02f2a: out <= 12'h72f;
      20'h02f2b: out <= 12'h72f;
      20'h02f2c: out <= 12'hfff;
      20'h02f2d: out <= 12'hc7f;
      20'h02f2e: out <= 12'hc7f;
      20'h02f2f: out <= 12'h72f;
      20'h02f30: out <= 12'h72f;
      20'h02f31: out <= 12'h72f;
      20'h02f32: out <= 12'hc7f;
      20'h02f33: out <= 12'hc7f;
      20'h02f34: out <= 12'hfff;
      20'h02f35: out <= 12'h72f;
      20'h02f36: out <= 12'h72f;
      20'h02f37: out <= 12'hc7f;
      20'h02f38: out <= 12'h000;
      20'h02f39: out <= 12'hc7f;
      20'h02f3a: out <= 12'hfff;
      20'h02f3b: out <= 12'h72f;
      20'h02f3c: out <= 12'hfff;
      20'h02f3d: out <= 12'hc7f;
      20'h02f3e: out <= 12'hc7f;
      20'h02f3f: out <= 12'h72f;
      20'h02f40: out <= 12'h72f;
      20'h02f41: out <= 12'h72f;
      20'h02f42: out <= 12'hc7f;
      20'h02f43: out <= 12'hc7f;
      20'h02f44: out <= 12'hfff;
      20'h02f45: out <= 12'h72f;
      20'h02f46: out <= 12'hfff;
      20'h02f47: out <= 12'hc7f;
      20'h02f48: out <= 12'h222;
      20'h02f49: out <= 12'h222;
      20'h02f4a: out <= 12'h222;
      20'h02f4b: out <= 12'h222;
      20'h02f4c: out <= 12'h222;
      20'h02f4d: out <= 12'h72f;
      20'h02f4e: out <= 12'hfff;
      20'h02f4f: out <= 12'hc7f;
      20'h02f50: out <= 12'hc7f;
      20'h02f51: out <= 12'hc7f;
      20'h02f52: out <= 12'hc7f;
      20'h02f53: out <= 12'hfff;
      20'h02f54: out <= 12'h72f;
      20'h02f55: out <= 12'h222;
      20'h02f56: out <= 12'h222;
      20'h02f57: out <= 12'h222;
      20'h02f58: out <= 12'h000;
      20'h02f59: out <= 12'h000;
      20'h02f5a: out <= 12'h000;
      20'h02f5b: out <= 12'h000;
      20'h02f5c: out <= 12'h000;
      20'h02f5d: out <= 12'h72f;
      20'h02f5e: out <= 12'hfff;
      20'h02f5f: out <= 12'hc7f;
      20'h02f60: out <= 12'hc7f;
      20'h02f61: out <= 12'hc7f;
      20'h02f62: out <= 12'hc7f;
      20'h02f63: out <= 12'hfff;
      20'h02f64: out <= 12'h72f;
      20'h02f65: out <= 12'h000;
      20'h02f66: out <= 12'h000;
      20'h02f67: out <= 12'h000;
      20'h02f68: out <= 12'h222;
      20'h02f69: out <= 12'hc7f;
      20'h02f6a: out <= 12'hfff;
      20'h02f6b: out <= 12'hc7f;
      20'h02f6c: out <= 12'h222;
      20'h02f6d: out <= 12'h72f;
      20'h02f6e: out <= 12'h72f;
      20'h02f6f: out <= 12'h72f;
      20'h02f70: out <= 12'hfff;
      20'h02f71: out <= 12'h72f;
      20'h02f72: out <= 12'h72f;
      20'h02f73: out <= 12'h72f;
      20'h02f74: out <= 12'h222;
      20'h02f75: out <= 12'hc7f;
      20'h02f76: out <= 12'hfff;
      20'h02f77: out <= 12'hc7f;
      20'h02f78: out <= 12'h000;
      20'h02f79: out <= 12'hc7f;
      20'h02f7a: out <= 12'h72f;
      20'h02f7b: out <= 12'hc7f;
      20'h02f7c: out <= 12'h000;
      20'h02f7d: out <= 12'h72f;
      20'h02f7e: out <= 12'h72f;
      20'h02f7f: out <= 12'h72f;
      20'h02f80: out <= 12'hfff;
      20'h02f81: out <= 12'h72f;
      20'h02f82: out <= 12'h72f;
      20'h02f83: out <= 12'h72f;
      20'h02f84: out <= 12'h000;
      20'h02f85: out <= 12'hc7f;
      20'h02f86: out <= 12'h72f;
      20'h02f87: out <= 12'hc7f;
      20'h02f88: out <= 12'h603;
      20'h02f89: out <= 12'h603;
      20'h02f8a: out <= 12'h603;
      20'h02f8b: out <= 12'h603;
      20'h02f8c: out <= 12'h6af;
      20'h02f8d: out <= 12'h4cd;
      20'h02f8e: out <= 12'h4cd;
      20'h02f8f: out <= 12'h6af;
      20'h02f90: out <= 12'hfff;
      20'h02f91: out <= 12'h4cd;
      20'h02f92: out <= 12'h4cd;
      20'h02f93: out <= 12'hfff;
      20'h02f94: out <= 12'h6af;
      20'h02f95: out <= 12'h4cd;
      20'h02f96: out <= 12'h4cd;
      20'h02f97: out <= 12'h6af;
      20'h02f98: out <= 12'hfff;
      20'h02f99: out <= 12'h4cd;
      20'h02f9a: out <= 12'h4cd;
      20'h02f9b: out <= 12'hfff;
      20'h02f9c: out <= 12'h380;
      20'h02f9d: out <= 12'hfff;
      20'h02f9e: out <= 12'h8d0;
      20'h02f9f: out <= 12'h8d0;
      20'h02fa0: out <= 12'h380;
      20'h02fa1: out <= 12'h000;
      20'h02fa2: out <= 12'h8d0;
      20'h02fa3: out <= 12'h000;
      20'h02fa4: out <= 12'h380;
      20'h02fa5: out <= 12'hfff;
      20'h02fa6: out <= 12'h8d0;
      20'h02fa7: out <= 12'h8d0;
      20'h02fa8: out <= 12'h380;
      20'h02fa9: out <= 12'h000;
      20'h02faa: out <= 12'h8d0;
      20'h02fab: out <= 12'h000;
      20'h02fac: out <= 12'h000;
      20'h02fad: out <= 12'h000;
      20'h02fae: out <= 12'hbbb;
      20'h02faf: out <= 12'hfff;
      20'h02fb0: out <= 12'h000;
      20'h02fb1: out <= 12'h000;
      20'h02fb2: out <= 12'hbbb;
      20'h02fb3: out <= 12'hfff;
      20'h02fb4: out <= 12'h000;
      20'h02fb5: out <= 12'h000;
      20'h02fb6: out <= 12'hbbb;
      20'h02fb7: out <= 12'hfff;
      20'h02fb8: out <= 12'h000;
      20'h02fb9: out <= 12'h000;
      20'h02fba: out <= 12'hbbb;
      20'h02fbb: out <= 12'hfff;
      20'h02fbc: out <= 12'h000;
      20'h02fbd: out <= 12'h6af;
      20'h02fbe: out <= 12'h000;
      20'h02fbf: out <= 12'hfff;
      20'h02fc0: out <= 12'hfff;
      20'h02fc1: out <= 12'h000;
      20'h02fc2: out <= 12'h6af;
      20'h02fc3: out <= 12'h4cd;
      20'h02fc4: out <= 12'hfff;
      20'h02fc5: out <= 12'h000;
      20'h02fc6: out <= 12'h6af;
      20'h02fc7: out <= 12'h000;
      20'h02fc8: out <= 12'hfff;
      20'h02fc9: out <= 12'h000;
      20'h02fca: out <= 12'h4cd;
      20'h02fcb: out <= 12'h6af;
      20'h02fcc: out <= 12'h000;
      20'h02fcd: out <= 12'h6af;
      20'h02fce: out <= 12'h000;
      20'h02fcf: out <= 12'hfff;
      20'h02fd0: out <= 12'h4cd;
      20'h02fd1: out <= 12'h000;
      20'h02fd2: out <= 12'h4cd;
      20'h02fd3: out <= 12'h000;
      20'h02fd4: out <= 12'h6af;
      20'h02fd5: out <= 12'h4cd;
      20'h02fd6: out <= 12'h4cd;
      20'h02fd7: out <= 12'hfff;
      20'h02fd8: out <= 12'hfff;
      20'h02fd9: out <= 12'h4cd;
      20'h02fda: out <= 12'h4cd;
      20'h02fdb: out <= 12'h000;
      20'h02fdc: out <= 12'h603;
      20'h02fdd: out <= 12'h603;
      20'h02fde: out <= 12'h603;
      20'h02fdf: out <= 12'h603;
      20'h02fe0: out <= 12'hee9;
      20'h02fe1: out <= 12'hf87;
      20'h02fe2: out <= 12'hee9;
      20'h02fe3: out <= 12'hf87;
      20'h02fe4: out <= 12'hf87;
      20'h02fe5: out <= 12'hb27;
      20'h02fe6: out <= 12'hf87;
      20'h02fe7: out <= 12'hb27;
      20'h02fe8: out <= 12'h000;
      20'h02fe9: out <= 12'h000;
      20'h02fea: out <= 12'h000;
      20'h02feb: out <= 12'h000;
      20'h02fec: out <= 12'h000;
      20'h02fed: out <= 12'h000;
      20'h02fee: out <= 12'h000;
      20'h02fef: out <= 12'h000;
      20'h02ff0: out <= 12'h000;
      20'h02ff1: out <= 12'h000;
      20'h02ff2: out <= 12'h000;
      20'h02ff3: out <= 12'h000;
      20'h02ff4: out <= 12'h000;
      20'h02ff5: out <= 12'h000;
      20'h02ff6: out <= 12'h000;
      20'h02ff7: out <= 12'h000;
      20'h02ff8: out <= 12'h916;
      20'h02ff9: out <= 12'h916;
      20'h02ffa: out <= 12'h916;
      20'h02ffb: out <= 12'h916;
      20'h02ffc: out <= 12'h916;
      20'h02ffd: out <= 12'h916;
      20'h02ffe: out <= 12'h916;
      20'h02fff: out <= 12'h916;
      20'h03000: out <= 12'hd29;
      20'h03001: out <= 12'hd29;
      20'h03002: out <= 12'hd29;
      20'h03003: out <= 12'hd29;
      20'h03004: out <= 12'hd29;
      20'h03005: out <= 12'hd29;
      20'h03006: out <= 12'hd29;
      20'h03007: out <= 12'hd29;
      20'h03008: out <= 12'h000;
      20'h03009: out <= 12'h000;
      20'h0300a: out <= 12'h000;
      20'h0300b: out <= 12'h000;
      20'h0300c: out <= 12'h000;
      20'h0300d: out <= 12'h000;
      20'h0300e: out <= 12'h000;
      20'h0300f: out <= 12'h000;
      20'h03010: out <= 12'h000;
      20'h03011: out <= 12'h000;
      20'h03012: out <= 12'h000;
      20'h03013: out <= 12'h000;
      20'h03014: out <= 12'h000;
      20'h03015: out <= 12'h000;
      20'h03016: out <= 12'h000;
      20'h03017: out <= 12'h000;
      20'h03018: out <= 12'h000;
      20'h03019: out <= 12'h000;
      20'h0301a: out <= 12'h000;
      20'h0301b: out <= 12'h000;
      20'h0301c: out <= 12'h000;
      20'h0301d: out <= 12'h000;
      20'h0301e: out <= 12'h000;
      20'h0301f: out <= 12'h000;
      20'h03020: out <= 12'h222;
      20'h03021: out <= 12'hc7f;
      20'h03022: out <= 12'hc7f;
      20'h03023: out <= 12'hc7f;
      20'h03024: out <= 12'h72f;
      20'h03025: out <= 12'h72f;
      20'h03026: out <= 12'h72f;
      20'h03027: out <= 12'h72f;
      20'h03028: out <= 12'h72f;
      20'h03029: out <= 12'h72f;
      20'h0302a: out <= 12'h72f;
      20'h0302b: out <= 12'hc7f;
      20'h0302c: out <= 12'hc7f;
      20'h0302d: out <= 12'h222;
      20'h0302e: out <= 12'h222;
      20'h0302f: out <= 12'h222;
      20'h03030: out <= 12'h000;
      20'h03031: out <= 12'hc7f;
      20'h03032: out <= 12'hc7f;
      20'h03033: out <= 12'hc7f;
      20'h03034: out <= 12'h72f;
      20'h03035: out <= 12'h72f;
      20'h03036: out <= 12'h72f;
      20'h03037: out <= 12'h72f;
      20'h03038: out <= 12'h72f;
      20'h03039: out <= 12'h72f;
      20'h0303a: out <= 12'h72f;
      20'h0303b: out <= 12'hc7f;
      20'h0303c: out <= 12'hc7f;
      20'h0303d: out <= 12'h000;
      20'h0303e: out <= 12'h000;
      20'h0303f: out <= 12'h000;
      20'h03040: out <= 12'h222;
      20'h03041: out <= 12'hc7f;
      20'h03042: out <= 12'hfff;
      20'h03043: out <= 12'hc7f;
      20'h03044: out <= 12'h72f;
      20'h03045: out <= 12'hfff;
      20'h03046: out <= 12'hc7f;
      20'h03047: out <= 12'hc7f;
      20'h03048: out <= 12'hc7f;
      20'h03049: out <= 12'hc7f;
      20'h0304a: out <= 12'hc7f;
      20'h0304b: out <= 12'hfff;
      20'h0304c: out <= 12'h72f;
      20'h0304d: out <= 12'hc7f;
      20'h0304e: out <= 12'hfff;
      20'h0304f: out <= 12'hc7f;
      20'h03050: out <= 12'h000;
      20'h03051: out <= 12'hc7f;
      20'h03052: out <= 12'h72f;
      20'h03053: out <= 12'hc7f;
      20'h03054: out <= 12'h72f;
      20'h03055: out <= 12'hfff;
      20'h03056: out <= 12'hc7f;
      20'h03057: out <= 12'hc7f;
      20'h03058: out <= 12'hc7f;
      20'h03059: out <= 12'hc7f;
      20'h0305a: out <= 12'hc7f;
      20'h0305b: out <= 12'hfff;
      20'h0305c: out <= 12'h72f;
      20'h0305d: out <= 12'hc7f;
      20'h0305e: out <= 12'h72f;
      20'h0305f: out <= 12'hc7f;
      20'h03060: out <= 12'h222;
      20'h03061: out <= 12'h222;
      20'h03062: out <= 12'h222;
      20'h03063: out <= 12'hc7f;
      20'h03064: out <= 12'hc7f;
      20'h03065: out <= 12'h72f;
      20'h03066: out <= 12'h72f;
      20'h03067: out <= 12'h72f;
      20'h03068: out <= 12'h72f;
      20'h03069: out <= 12'h72f;
      20'h0306a: out <= 12'h72f;
      20'h0306b: out <= 12'h72f;
      20'h0306c: out <= 12'hc7f;
      20'h0306d: out <= 12'hc7f;
      20'h0306e: out <= 12'hc7f;
      20'h0306f: out <= 12'h222;
      20'h03070: out <= 12'h000;
      20'h03071: out <= 12'h000;
      20'h03072: out <= 12'h000;
      20'h03073: out <= 12'hc7f;
      20'h03074: out <= 12'hc7f;
      20'h03075: out <= 12'h72f;
      20'h03076: out <= 12'h72f;
      20'h03077: out <= 12'h72f;
      20'h03078: out <= 12'h72f;
      20'h03079: out <= 12'h72f;
      20'h0307a: out <= 12'h72f;
      20'h0307b: out <= 12'h72f;
      20'h0307c: out <= 12'hc7f;
      20'h0307d: out <= 12'hc7f;
      20'h0307e: out <= 12'hc7f;
      20'h0307f: out <= 12'h000;
      20'h03080: out <= 12'h222;
      20'h03081: out <= 12'hc7f;
      20'h03082: out <= 12'h72f;
      20'h03083: out <= 12'hc7f;
      20'h03084: out <= 12'h222;
      20'h03085: out <= 12'h222;
      20'h03086: out <= 12'h222;
      20'h03087: out <= 12'h72f;
      20'h03088: out <= 12'hfff;
      20'h03089: out <= 12'h72f;
      20'h0308a: out <= 12'h222;
      20'h0308b: out <= 12'h222;
      20'h0308c: out <= 12'h222;
      20'h0308d: out <= 12'hc7f;
      20'h0308e: out <= 12'h72f;
      20'h0308f: out <= 12'hc7f;
      20'h03090: out <= 12'h000;
      20'h03091: out <= 12'hc7f;
      20'h03092: out <= 12'hfff;
      20'h03093: out <= 12'hc7f;
      20'h03094: out <= 12'h000;
      20'h03095: out <= 12'h000;
      20'h03096: out <= 12'h000;
      20'h03097: out <= 12'h72f;
      20'h03098: out <= 12'hfff;
      20'h03099: out <= 12'h72f;
      20'h0309a: out <= 12'h000;
      20'h0309b: out <= 12'h000;
      20'h0309c: out <= 12'h000;
      20'h0309d: out <= 12'hc7f;
      20'h0309e: out <= 12'hfff;
      20'h0309f: out <= 12'hc7f;
      20'h030a0: out <= 12'h603;
      20'h030a1: out <= 12'h603;
      20'h030a2: out <= 12'h603;
      20'h030a3: out <= 12'h603;
      20'h030a4: out <= 12'hfff;
      20'h030a5: out <= 12'h6af;
      20'h030a6: out <= 12'h6af;
      20'h030a7: out <= 12'hfff;
      20'h030a8: out <= 12'h4cd;
      20'h030a9: out <= 12'h4cd;
      20'h030aa: out <= 12'h4cd;
      20'h030ab: out <= 12'h4cd;
      20'h030ac: out <= 12'hfff;
      20'h030ad: out <= 12'h6af;
      20'h030ae: out <= 12'h6af;
      20'h030af: out <= 12'hfff;
      20'h030b0: out <= 12'h4cd;
      20'h030b1: out <= 12'h4cd;
      20'h030b2: out <= 12'h4cd;
      20'h030b3: out <= 12'h4cd;
      20'h030b4: out <= 12'hfff;
      20'h030b5: out <= 12'h8d0;
      20'h030b6: out <= 12'h8d0;
      20'h030b7: out <= 12'h380;
      20'h030b8: out <= 12'h8d0;
      20'h030b9: out <= 12'h8d0;
      20'h030ba: out <= 12'h000;
      20'h030bb: out <= 12'h380;
      20'h030bc: out <= 12'hfff;
      20'h030bd: out <= 12'h8d0;
      20'h030be: out <= 12'h8d0;
      20'h030bf: out <= 12'h380;
      20'h030c0: out <= 12'h8d0;
      20'h030c1: out <= 12'h8d0;
      20'h030c2: out <= 12'h000;
      20'h030c3: out <= 12'h380;
      20'h030c4: out <= 12'hfff;
      20'h030c5: out <= 12'h666;
      20'h030c6: out <= 12'h000;
      20'h030c7: out <= 12'h000;
      20'h030c8: out <= 12'hfff;
      20'h030c9: out <= 12'h666;
      20'h030ca: out <= 12'h000;
      20'h030cb: out <= 12'h000;
      20'h030cc: out <= 12'hfff;
      20'h030cd: out <= 12'h666;
      20'h030ce: out <= 12'h000;
      20'h030cf: out <= 12'h000;
      20'h030d0: out <= 12'hfff;
      20'h030d1: out <= 12'h666;
      20'h030d2: out <= 12'h000;
      20'h030d3: out <= 12'h000;
      20'h030d4: out <= 12'h000;
      20'h030d5: out <= 12'h6af;
      20'h030d6: out <= 12'h000;
      20'h030d7: out <= 12'hfff;
      20'h030d8: out <= 12'hfff;
      20'h030d9: out <= 12'h000;
      20'h030da: out <= 12'h6af;
      20'h030db: out <= 12'h4cd;
      20'h030dc: out <= 12'hfff;
      20'h030dd: out <= 12'h000;
      20'h030de: out <= 12'h6af;
      20'h030df: out <= 12'h4cd;
      20'h030e0: out <= 12'hfff;
      20'h030e1: out <= 12'hfff;
      20'h030e2: out <= 12'h4cd;
      20'h030e3: out <= 12'h6af;
      20'h030e4: out <= 12'h000;
      20'h030e5: out <= 12'h6af;
      20'h030e6: out <= 12'h4cd;
      20'h030e7: out <= 12'hfff;
      20'h030e8: out <= 12'h4cd;
      20'h030e9: out <= 12'h000;
      20'h030ea: out <= 12'h000;
      20'h030eb: out <= 12'h000;
      20'h030ec: out <= 12'h6af;
      20'h030ed: out <= 12'hfff;
      20'h030ee: out <= 12'hfff;
      20'h030ef: out <= 12'h000;
      20'h030f0: out <= 12'hfff;
      20'h030f1: out <= 12'h4cd;
      20'h030f2: out <= 12'hfff;
      20'h030f3: out <= 12'h000;
      20'h030f4: out <= 12'h603;
      20'h030f5: out <= 12'h603;
      20'h030f6: out <= 12'h603;
      20'h030f7: out <= 12'h603;
      20'h030f8: out <= 12'hee9;
      20'h030f9: out <= 12'hf87;
      20'h030fa: out <= 12'hee9;
      20'h030fb: out <= 12'hf87;
      20'h030fc: out <= 12'hf87;
      20'h030fd: out <= 12'hb27;
      20'h030fe: out <= 12'hf87;
      20'h030ff: out <= 12'hb27;
      20'h03100: out <= 12'h000;
      20'h03101: out <= 12'h000;
      20'h03102: out <= 12'h000;
      20'h03103: out <= 12'h000;
      20'h03104: out <= 12'h000;
      20'h03105: out <= 12'h000;
      20'h03106: out <= 12'h000;
      20'h03107: out <= 12'h000;
      20'h03108: out <= 12'h000;
      20'h03109: out <= 12'h000;
      20'h0310a: out <= 12'h000;
      20'h0310b: out <= 12'h000;
      20'h0310c: out <= 12'h000;
      20'h0310d: out <= 12'h000;
      20'h0310e: out <= 12'h000;
      20'h0310f: out <= 12'h000;
      20'h03110: out <= 12'h916;
      20'h03111: out <= 12'h916;
      20'h03112: out <= 12'h916;
      20'h03113: out <= 12'h916;
      20'h03114: out <= 12'h916;
      20'h03115: out <= 12'h916;
      20'h03116: out <= 12'h916;
      20'h03117: out <= 12'h916;
      20'h03118: out <= 12'hd29;
      20'h03119: out <= 12'hd29;
      20'h0311a: out <= 12'hd29;
      20'h0311b: out <= 12'hd29;
      20'h0311c: out <= 12'hd29;
      20'h0311d: out <= 12'hd29;
      20'h0311e: out <= 12'hd29;
      20'h0311f: out <= 12'hd29;
      20'h03120: out <= 12'h000;
      20'h03121: out <= 12'h000;
      20'h03122: out <= 12'h000;
      20'h03123: out <= 12'h000;
      20'h03124: out <= 12'h000;
      20'h03125: out <= 12'h000;
      20'h03126: out <= 12'h000;
      20'h03127: out <= 12'h000;
      20'h03128: out <= 12'h000;
      20'h03129: out <= 12'h000;
      20'h0312a: out <= 12'h000;
      20'h0312b: out <= 12'h000;
      20'h0312c: out <= 12'h000;
      20'h0312d: out <= 12'h000;
      20'h0312e: out <= 12'h000;
      20'h0312f: out <= 12'h000;
      20'h03130: out <= 12'h000;
      20'h03131: out <= 12'h000;
      20'h03132: out <= 12'h000;
      20'h03133: out <= 12'h000;
      20'h03134: out <= 12'h000;
      20'h03135: out <= 12'h000;
      20'h03136: out <= 12'h000;
      20'h03137: out <= 12'h000;
      20'h03138: out <= 12'h222;
      20'h03139: out <= 12'hfff;
      20'h0313a: out <= 12'h72f;
      20'h0313b: out <= 12'hfff;
      20'h0313c: out <= 12'h72f;
      20'h0313d: out <= 12'hfff;
      20'h0313e: out <= 12'h72f;
      20'h0313f: out <= 12'hfff;
      20'h03140: out <= 12'h72f;
      20'h03141: out <= 12'hfff;
      20'h03142: out <= 12'h72f;
      20'h03143: out <= 12'hfff;
      20'h03144: out <= 12'h72f;
      20'h03145: out <= 12'h222;
      20'h03146: out <= 12'h222;
      20'h03147: out <= 12'h222;
      20'h03148: out <= 12'h000;
      20'h03149: out <= 12'hc7f;
      20'h0314a: out <= 12'hfff;
      20'h0314b: out <= 12'h72f;
      20'h0314c: out <= 12'hfff;
      20'h0314d: out <= 12'h72f;
      20'h0314e: out <= 12'hfff;
      20'h0314f: out <= 12'h72f;
      20'h03150: out <= 12'hfff;
      20'h03151: out <= 12'h72f;
      20'h03152: out <= 12'hfff;
      20'h03153: out <= 12'h72f;
      20'h03154: out <= 12'hfff;
      20'h03155: out <= 12'h000;
      20'h03156: out <= 12'h000;
      20'h03157: out <= 12'h000;
      20'h03158: out <= 12'h222;
      20'h03159: out <= 12'hc7f;
      20'h0315a: out <= 12'h72f;
      20'h0315b: out <= 12'hc7f;
      20'h0315c: out <= 12'h222;
      20'h0315d: out <= 12'h72f;
      20'h0315e: out <= 12'h72f;
      20'h0315f: out <= 12'h72f;
      20'h03160: out <= 12'h72f;
      20'h03161: out <= 12'h72f;
      20'h03162: out <= 12'h72f;
      20'h03163: out <= 12'h72f;
      20'h03164: out <= 12'h222;
      20'h03165: out <= 12'hc7f;
      20'h03166: out <= 12'h72f;
      20'h03167: out <= 12'hc7f;
      20'h03168: out <= 12'h000;
      20'h03169: out <= 12'hc7f;
      20'h0316a: out <= 12'hfff;
      20'h0316b: out <= 12'hc7f;
      20'h0316c: out <= 12'h000;
      20'h0316d: out <= 12'h72f;
      20'h0316e: out <= 12'h72f;
      20'h0316f: out <= 12'h72f;
      20'h03170: out <= 12'h72f;
      20'h03171: out <= 12'h72f;
      20'h03172: out <= 12'h72f;
      20'h03173: out <= 12'h72f;
      20'h03174: out <= 12'h000;
      20'h03175: out <= 12'hc7f;
      20'h03176: out <= 12'hfff;
      20'h03177: out <= 12'hc7f;
      20'h03178: out <= 12'h222;
      20'h03179: out <= 12'h222;
      20'h0317a: out <= 12'h222;
      20'h0317b: out <= 12'h72f;
      20'h0317c: out <= 12'hfff;
      20'h0317d: out <= 12'h72f;
      20'h0317e: out <= 12'hfff;
      20'h0317f: out <= 12'h72f;
      20'h03180: out <= 12'hfff;
      20'h03181: out <= 12'h72f;
      20'h03182: out <= 12'hfff;
      20'h03183: out <= 12'h72f;
      20'h03184: out <= 12'hfff;
      20'h03185: out <= 12'h72f;
      20'h03186: out <= 12'hfff;
      20'h03187: out <= 12'h222;
      20'h03188: out <= 12'h000;
      20'h03189: out <= 12'h000;
      20'h0318a: out <= 12'h000;
      20'h0318b: out <= 12'hfff;
      20'h0318c: out <= 12'h72f;
      20'h0318d: out <= 12'hfff;
      20'h0318e: out <= 12'h72f;
      20'h0318f: out <= 12'hfff;
      20'h03190: out <= 12'h72f;
      20'h03191: out <= 12'hfff;
      20'h03192: out <= 12'h72f;
      20'h03193: out <= 12'hfff;
      20'h03194: out <= 12'h72f;
      20'h03195: out <= 12'hfff;
      20'h03196: out <= 12'hc7f;
      20'h03197: out <= 12'h000;
      20'h03198: out <= 12'h222;
      20'h03199: out <= 12'h222;
      20'h0319a: out <= 12'h222;
      20'h0319b: out <= 12'h222;
      20'h0319c: out <= 12'h222;
      20'h0319d: out <= 12'h222;
      20'h0319e: out <= 12'h222;
      20'h0319f: out <= 12'h72f;
      20'h031a0: out <= 12'hfff;
      20'h031a1: out <= 12'h72f;
      20'h031a2: out <= 12'h222;
      20'h031a3: out <= 12'h222;
      20'h031a4: out <= 12'h222;
      20'h031a5: out <= 12'h222;
      20'h031a6: out <= 12'h222;
      20'h031a7: out <= 12'h222;
      20'h031a8: out <= 12'h000;
      20'h031a9: out <= 12'h000;
      20'h031aa: out <= 12'h000;
      20'h031ab: out <= 12'h000;
      20'h031ac: out <= 12'h000;
      20'h031ad: out <= 12'h000;
      20'h031ae: out <= 12'h000;
      20'h031af: out <= 12'h72f;
      20'h031b0: out <= 12'hfff;
      20'h031b1: out <= 12'h72f;
      20'h031b2: out <= 12'h000;
      20'h031b3: out <= 12'h000;
      20'h031b4: out <= 12'h000;
      20'h031b5: out <= 12'h000;
      20'h031b6: out <= 12'h000;
      20'h031b7: out <= 12'h000;
      20'h031b8: out <= 12'h603;
      20'h031b9: out <= 12'h603;
      20'h031ba: out <= 12'h603;
      20'h031bb: out <= 12'h603;
      20'h031bc: out <= 12'h4cd;
      20'h031bd: out <= 12'hfff;
      20'h031be: out <= 12'hfff;
      20'h031bf: out <= 12'h4cd;
      20'h031c0: out <= 12'h4cd;
      20'h031c1: out <= 12'h6af;
      20'h031c2: out <= 12'h6af;
      20'h031c3: out <= 12'h4cd;
      20'h031c4: out <= 12'h4cd;
      20'h031c5: out <= 12'hfff;
      20'h031c6: out <= 12'hfff;
      20'h031c7: out <= 12'h4cd;
      20'h031c8: out <= 12'h4cd;
      20'h031c9: out <= 12'h6af;
      20'h031ca: out <= 12'h6af;
      20'h031cb: out <= 12'h4cd;
      20'h031cc: out <= 12'h380;
      20'h031cd: out <= 12'h8d0;
      20'h031ce: out <= 12'h380;
      20'h031cf: out <= 12'h380;
      20'h031d0: out <= 12'h8d0;
      20'h031d1: out <= 12'h380;
      20'h031d2: out <= 12'h380;
      20'h031d3: out <= 12'h380;
      20'h031d4: out <= 12'h380;
      20'h031d5: out <= 12'h8d0;
      20'h031d6: out <= 12'h380;
      20'h031d7: out <= 12'h380;
      20'h031d8: out <= 12'h8d0;
      20'h031d9: out <= 12'h380;
      20'h031da: out <= 12'h380;
      20'h031db: out <= 12'h380;
      20'h031dc: out <= 12'hbbb;
      20'h031dd: out <= 12'hfff;
      20'h031de: out <= 12'h000;
      20'h031df: out <= 12'h000;
      20'h031e0: out <= 12'hbbb;
      20'h031e1: out <= 12'hfff;
      20'h031e2: out <= 12'h000;
      20'h031e3: out <= 12'h000;
      20'h031e4: out <= 12'hbbb;
      20'h031e5: out <= 12'hfff;
      20'h031e6: out <= 12'h000;
      20'h031e7: out <= 12'h000;
      20'h031e8: out <= 12'hbbb;
      20'h031e9: out <= 12'hfff;
      20'h031ea: out <= 12'h000;
      20'h031eb: out <= 12'h000;
      20'h031ec: out <= 12'h000;
      20'h031ed: out <= 12'h6af;
      20'h031ee: out <= 12'h4cd;
      20'h031ef: out <= 12'hfff;
      20'h031f0: out <= 12'hfff;
      20'h031f1: out <= 12'h000;
      20'h031f2: out <= 12'h6af;
      20'h031f3: out <= 12'h4cd;
      20'h031f4: out <= 12'hfff;
      20'h031f5: out <= 12'h000;
      20'h031f6: out <= 12'h6af;
      20'h031f7: out <= 12'h4cd;
      20'h031f8: out <= 12'hfff;
      20'h031f9: out <= 12'hfff;
      20'h031fa: out <= 12'h4cd;
      20'h031fb: out <= 12'h6af;
      20'h031fc: out <= 12'h000;
      20'h031fd: out <= 12'h6af;
      20'h031fe: out <= 12'h4cd;
      20'h031ff: out <= 12'hfff;
      20'h03200: out <= 12'h4cd;
      20'h03201: out <= 12'h000;
      20'h03202: out <= 12'h6af;
      20'h03203: out <= 12'h4cd;
      20'h03204: out <= 12'h4cd;
      20'h03205: out <= 12'h4cd;
      20'h03206: out <= 12'hfff;
      20'h03207: out <= 12'hfff;
      20'h03208: out <= 12'hfff;
      20'h03209: out <= 12'h000;
      20'h0320a: out <= 12'h000;
      20'h0320b: out <= 12'h6af;
      20'h0320c: out <= 12'h603;
      20'h0320d: out <= 12'h603;
      20'h0320e: out <= 12'h603;
      20'h0320f: out <= 12'h603;
      20'h03210: out <= 12'hee9;
      20'h03211: out <= 12'hf87;
      20'h03212: out <= 12'hee9;
      20'h03213: out <= 12'hb27;
      20'h03214: out <= 12'hb27;
      20'h03215: out <= 12'hb27;
      20'h03216: out <= 12'hf87;
      20'h03217: out <= 12'hb27;
      20'h03218: out <= 12'h000;
      20'h03219: out <= 12'h000;
      20'h0321a: out <= 12'h000;
      20'h0321b: out <= 12'h000;
      20'h0321c: out <= 12'h000;
      20'h0321d: out <= 12'h000;
      20'h0321e: out <= 12'h000;
      20'h0321f: out <= 12'h000;
      20'h03220: out <= 12'h000;
      20'h03221: out <= 12'h000;
      20'h03222: out <= 12'h000;
      20'h03223: out <= 12'h000;
      20'h03224: out <= 12'h000;
      20'h03225: out <= 12'h000;
      20'h03226: out <= 12'h000;
      20'h03227: out <= 12'h000;
      20'h03228: out <= 12'h916;
      20'h03229: out <= 12'h916;
      20'h0322a: out <= 12'h916;
      20'h0322b: out <= 12'h916;
      20'h0322c: out <= 12'h916;
      20'h0322d: out <= 12'h916;
      20'h0322e: out <= 12'h916;
      20'h0322f: out <= 12'h916;
      20'h03230: out <= 12'hd29;
      20'h03231: out <= 12'hd29;
      20'h03232: out <= 12'hd29;
      20'h03233: out <= 12'hd29;
      20'h03234: out <= 12'hd29;
      20'h03235: out <= 12'hd29;
      20'h03236: out <= 12'hd29;
      20'h03237: out <= 12'hd29;
      20'h03238: out <= 12'h000;
      20'h03239: out <= 12'h000;
      20'h0323a: out <= 12'h000;
      20'h0323b: out <= 12'h000;
      20'h0323c: out <= 12'h000;
      20'h0323d: out <= 12'h000;
      20'h0323e: out <= 12'h000;
      20'h0323f: out <= 12'h000;
      20'h03240: out <= 12'h000;
      20'h03241: out <= 12'h000;
      20'h03242: out <= 12'h000;
      20'h03243: out <= 12'h000;
      20'h03244: out <= 12'h000;
      20'h03245: out <= 12'h000;
      20'h03246: out <= 12'h000;
      20'h03247: out <= 12'h000;
      20'h03248: out <= 12'h000;
      20'h03249: out <= 12'h000;
      20'h0324a: out <= 12'h000;
      20'h0324b: out <= 12'h000;
      20'h0324c: out <= 12'h000;
      20'h0324d: out <= 12'h000;
      20'h0324e: out <= 12'h000;
      20'h0324f: out <= 12'h000;
      20'h03250: out <= 12'h222;
      20'h03251: out <= 12'hc7f;
      20'h03252: out <= 12'hc7f;
      20'h03253: out <= 12'hc7f;
      20'h03254: out <= 12'hc7f;
      20'h03255: out <= 12'hc7f;
      20'h03256: out <= 12'hc7f;
      20'h03257: out <= 12'hc7f;
      20'h03258: out <= 12'hc7f;
      20'h03259: out <= 12'hc7f;
      20'h0325a: out <= 12'hc7f;
      20'h0325b: out <= 12'hc7f;
      20'h0325c: out <= 12'hc7f;
      20'h0325d: out <= 12'h222;
      20'h0325e: out <= 12'h222;
      20'h0325f: out <= 12'h222;
      20'h03260: out <= 12'h000;
      20'h03261: out <= 12'hc7f;
      20'h03262: out <= 12'hc7f;
      20'h03263: out <= 12'hc7f;
      20'h03264: out <= 12'hc7f;
      20'h03265: out <= 12'hc7f;
      20'h03266: out <= 12'hc7f;
      20'h03267: out <= 12'hc7f;
      20'h03268: out <= 12'hc7f;
      20'h03269: out <= 12'hc7f;
      20'h0326a: out <= 12'hc7f;
      20'h0326b: out <= 12'hc7f;
      20'h0326c: out <= 12'hc7f;
      20'h0326d: out <= 12'h000;
      20'h0326e: out <= 12'h000;
      20'h0326f: out <= 12'h000;
      20'h03270: out <= 12'h222;
      20'h03271: out <= 12'hc7f;
      20'h03272: out <= 12'hfff;
      20'h03273: out <= 12'hc7f;
      20'h03274: out <= 12'h222;
      20'h03275: out <= 12'h222;
      20'h03276: out <= 12'h222;
      20'h03277: out <= 12'h222;
      20'h03278: out <= 12'h222;
      20'h03279: out <= 12'h222;
      20'h0327a: out <= 12'h222;
      20'h0327b: out <= 12'h222;
      20'h0327c: out <= 12'h222;
      20'h0327d: out <= 12'hc7f;
      20'h0327e: out <= 12'hfff;
      20'h0327f: out <= 12'hc7f;
      20'h03280: out <= 12'h000;
      20'h03281: out <= 12'hc7f;
      20'h03282: out <= 12'hc7f;
      20'h03283: out <= 12'hc7f;
      20'h03284: out <= 12'h000;
      20'h03285: out <= 12'h000;
      20'h03286: out <= 12'h000;
      20'h03287: out <= 12'h000;
      20'h03288: out <= 12'h000;
      20'h03289: out <= 12'h000;
      20'h0328a: out <= 12'h000;
      20'h0328b: out <= 12'h000;
      20'h0328c: out <= 12'h000;
      20'h0328d: out <= 12'hc7f;
      20'h0328e: out <= 12'hc7f;
      20'h0328f: out <= 12'hc7f;
      20'h03290: out <= 12'h222;
      20'h03291: out <= 12'h222;
      20'h03292: out <= 12'h222;
      20'h03293: out <= 12'hc7f;
      20'h03294: out <= 12'hc7f;
      20'h03295: out <= 12'hc7f;
      20'h03296: out <= 12'hc7f;
      20'h03297: out <= 12'hc7f;
      20'h03298: out <= 12'hc7f;
      20'h03299: out <= 12'hc7f;
      20'h0329a: out <= 12'hc7f;
      20'h0329b: out <= 12'hc7f;
      20'h0329c: out <= 12'hc7f;
      20'h0329d: out <= 12'hc7f;
      20'h0329e: out <= 12'hc7f;
      20'h0329f: out <= 12'h222;
      20'h032a0: out <= 12'h000;
      20'h032a1: out <= 12'h000;
      20'h032a2: out <= 12'h000;
      20'h032a3: out <= 12'hc7f;
      20'h032a4: out <= 12'hc7f;
      20'h032a5: out <= 12'hc7f;
      20'h032a6: out <= 12'hc7f;
      20'h032a7: out <= 12'hc7f;
      20'h032a8: out <= 12'hc7f;
      20'h032a9: out <= 12'hc7f;
      20'h032aa: out <= 12'hc7f;
      20'h032ab: out <= 12'hc7f;
      20'h032ac: out <= 12'hc7f;
      20'h032ad: out <= 12'hc7f;
      20'h032ae: out <= 12'hc7f;
      20'h032af: out <= 12'h000;
      20'h032b0: out <= 12'h222;
      20'h032b1: out <= 12'h222;
      20'h032b2: out <= 12'h222;
      20'h032b3: out <= 12'h222;
      20'h032b4: out <= 12'h222;
      20'h032b5: out <= 12'h222;
      20'h032b6: out <= 12'h222;
      20'h032b7: out <= 12'h72f;
      20'h032b8: out <= 12'hfff;
      20'h032b9: out <= 12'h72f;
      20'h032ba: out <= 12'h222;
      20'h032bb: out <= 12'h222;
      20'h032bc: out <= 12'h222;
      20'h032bd: out <= 12'h222;
      20'h032be: out <= 12'h222;
      20'h032bf: out <= 12'h222;
      20'h032c0: out <= 12'h000;
      20'h032c1: out <= 12'h000;
      20'h032c2: out <= 12'h000;
      20'h032c3: out <= 12'h000;
      20'h032c4: out <= 12'h000;
      20'h032c5: out <= 12'h000;
      20'h032c6: out <= 12'h000;
      20'h032c7: out <= 12'h72f;
      20'h032c8: out <= 12'hfff;
      20'h032c9: out <= 12'h72f;
      20'h032ca: out <= 12'h000;
      20'h032cb: out <= 12'h000;
      20'h032cc: out <= 12'h000;
      20'h032cd: out <= 12'h000;
      20'h032ce: out <= 12'h000;
      20'h032cf: out <= 12'h000;
      20'h032d0: out <= 12'h603;
      20'h032d1: out <= 12'h603;
      20'h032d2: out <= 12'h603;
      20'h032d3: out <= 12'h603;
      20'h032d4: out <= 12'h4cd;
      20'h032d5: out <= 12'h4cd;
      20'h032d6: out <= 12'h4cd;
      20'h032d7: out <= 12'h4cd;
      20'h032d8: out <= 12'h6af;
      20'h032d9: out <= 12'hfff;
      20'h032da: out <= 12'hfff;
      20'h032db: out <= 12'h6af;
      20'h032dc: out <= 12'h4cd;
      20'h032dd: out <= 12'h4cd;
      20'h032de: out <= 12'h4cd;
      20'h032df: out <= 12'h4cd;
      20'h032e0: out <= 12'h6af;
      20'h032e1: out <= 12'hfff;
      20'h032e2: out <= 12'hfff;
      20'h032e3: out <= 12'h6af;
      20'h032e4: out <= 12'h000;
      20'h032e5: out <= 12'h380;
      20'h032e6: out <= 12'h8d0;
      20'h032e7: out <= 12'h8d0;
      20'h032e8: out <= 12'h000;
      20'h032e9: out <= 12'h380;
      20'h032ea: out <= 12'h000;
      20'h032eb: out <= 12'h380;
      20'h032ec: out <= 12'h000;
      20'h032ed: out <= 12'h380;
      20'h032ee: out <= 12'h8d0;
      20'h032ef: out <= 12'h8d0;
      20'h032f0: out <= 12'h000;
      20'h032f1: out <= 12'h380;
      20'h032f2: out <= 12'h000;
      20'h032f3: out <= 12'h380;
      20'h032f4: out <= 12'h000;
      20'h032f5: out <= 12'h000;
      20'h032f6: out <= 12'hfff;
      20'h032f7: out <= 12'h666;
      20'h032f8: out <= 12'h000;
      20'h032f9: out <= 12'h000;
      20'h032fa: out <= 12'hfff;
      20'h032fb: out <= 12'h666;
      20'h032fc: out <= 12'h000;
      20'h032fd: out <= 12'h000;
      20'h032fe: out <= 12'hfff;
      20'h032ff: out <= 12'h666;
      20'h03300: out <= 12'h000;
      20'h03301: out <= 12'h000;
      20'h03302: out <= 12'hfff;
      20'h03303: out <= 12'h666;
      20'h03304: out <= 12'h000;
      20'h03305: out <= 12'h000;
      20'h03306: out <= 12'h000;
      20'h03307: out <= 12'h000;
      20'h03308: out <= 12'h000;
      20'h03309: out <= 12'h000;
      20'h0330a: out <= 12'h000;
      20'h0330b: out <= 12'h000;
      20'h0330c: out <= 12'h000;
      20'h0330d: out <= 12'h000;
      20'h0330e: out <= 12'h000;
      20'h0330f: out <= 12'h000;
      20'h03310: out <= 12'h000;
      20'h03311: out <= 12'h000;
      20'h03312: out <= 12'h000;
      20'h03313: out <= 12'h000;
      20'h03314: out <= 12'h000;
      20'h03315: out <= 12'h000;
      20'h03316: out <= 12'h000;
      20'h03317: out <= 12'h000;
      20'h03318: out <= 12'h000;
      20'h03319: out <= 12'h000;
      20'h0331a: out <= 12'h000;
      20'h0331b: out <= 12'h000;
      20'h0331c: out <= 12'h000;
      20'h0331d: out <= 12'h000;
      20'h0331e: out <= 12'h000;
      20'h0331f: out <= 12'h000;
      20'h03320: out <= 12'h000;
      20'h03321: out <= 12'h000;
      20'h03322: out <= 12'h000;
      20'h03323: out <= 12'h000;
      20'h03324: out <= 12'h603;
      20'h03325: out <= 12'h603;
      20'h03326: out <= 12'h603;
      20'h03327: out <= 12'h603;
      20'h03328: out <= 12'hee9;
      20'h03329: out <= 12'hf87;
      20'h0332a: out <= 12'hf87;
      20'h0332b: out <= 12'hf87;
      20'h0332c: out <= 12'hf87;
      20'h0332d: out <= 12'hf87;
      20'h0332e: out <= 12'hf87;
      20'h0332f: out <= 12'hb27;
      20'h03330: out <= 12'h000;
      20'h03331: out <= 12'h000;
      20'h03332: out <= 12'h000;
      20'h03333: out <= 12'h000;
      20'h03334: out <= 12'h000;
      20'h03335: out <= 12'h000;
      20'h03336: out <= 12'h000;
      20'h03337: out <= 12'h000;
      20'h03338: out <= 12'h000;
      20'h03339: out <= 12'h000;
      20'h0333a: out <= 12'h000;
      20'h0333b: out <= 12'h000;
      20'h0333c: out <= 12'h000;
      20'h0333d: out <= 12'h000;
      20'h0333e: out <= 12'h000;
      20'h0333f: out <= 12'h000;
      20'h03340: out <= 12'h916;
      20'h03341: out <= 12'h916;
      20'h03342: out <= 12'h916;
      20'h03343: out <= 12'h916;
      20'h03344: out <= 12'h916;
      20'h03345: out <= 12'h916;
      20'h03346: out <= 12'h916;
      20'h03347: out <= 12'h916;
      20'h03348: out <= 12'hd29;
      20'h03349: out <= 12'hd29;
      20'h0334a: out <= 12'hd29;
      20'h0334b: out <= 12'hd29;
      20'h0334c: out <= 12'hd29;
      20'h0334d: out <= 12'hd29;
      20'h0334e: out <= 12'hd29;
      20'h0334f: out <= 12'hd29;
      20'h03350: out <= 12'h000;
      20'h03351: out <= 12'h000;
      20'h03352: out <= 12'h000;
      20'h03353: out <= 12'h000;
      20'h03354: out <= 12'h000;
      20'h03355: out <= 12'h000;
      20'h03356: out <= 12'h000;
      20'h03357: out <= 12'h000;
      20'h03358: out <= 12'h000;
      20'h03359: out <= 12'h000;
      20'h0335a: out <= 12'h000;
      20'h0335b: out <= 12'h000;
      20'h0335c: out <= 12'h000;
      20'h0335d: out <= 12'h000;
      20'h0335e: out <= 12'h000;
      20'h0335f: out <= 12'h000;
      20'h03360: out <= 12'h000;
      20'h03361: out <= 12'h000;
      20'h03362: out <= 12'h000;
      20'h03363: out <= 12'h000;
      20'h03364: out <= 12'h000;
      20'h03365: out <= 12'h000;
      20'h03366: out <= 12'h000;
      20'h03367: out <= 12'h000;
      20'h03368: out <= 12'h222;
      20'h03369: out <= 12'h222;
      20'h0336a: out <= 12'h222;
      20'h0336b: out <= 12'h222;
      20'h0336c: out <= 12'h222;
      20'h0336d: out <= 12'h222;
      20'h0336e: out <= 12'h222;
      20'h0336f: out <= 12'h222;
      20'h03370: out <= 12'h222;
      20'h03371: out <= 12'h222;
      20'h03372: out <= 12'h222;
      20'h03373: out <= 12'h222;
      20'h03374: out <= 12'h222;
      20'h03375: out <= 12'h222;
      20'h03376: out <= 12'h222;
      20'h03377: out <= 12'h222;
      20'h03378: out <= 12'h000;
      20'h03379: out <= 12'h000;
      20'h0337a: out <= 12'h000;
      20'h0337b: out <= 12'h000;
      20'h0337c: out <= 12'h000;
      20'h0337d: out <= 12'h000;
      20'h0337e: out <= 12'h000;
      20'h0337f: out <= 12'h000;
      20'h03380: out <= 12'h000;
      20'h03381: out <= 12'h000;
      20'h03382: out <= 12'h000;
      20'h03383: out <= 12'h000;
      20'h03384: out <= 12'h000;
      20'h03385: out <= 12'h000;
      20'h03386: out <= 12'h000;
      20'h03387: out <= 12'h000;
      20'h03388: out <= 12'h222;
      20'h03389: out <= 12'h222;
      20'h0338a: out <= 12'h222;
      20'h0338b: out <= 12'h222;
      20'h0338c: out <= 12'h222;
      20'h0338d: out <= 12'h222;
      20'h0338e: out <= 12'h222;
      20'h0338f: out <= 12'h222;
      20'h03390: out <= 12'h222;
      20'h03391: out <= 12'h222;
      20'h03392: out <= 12'h222;
      20'h03393: out <= 12'h222;
      20'h03394: out <= 12'h222;
      20'h03395: out <= 12'h222;
      20'h03396: out <= 12'h222;
      20'h03397: out <= 12'h222;
      20'h03398: out <= 12'h000;
      20'h03399: out <= 12'h000;
      20'h0339a: out <= 12'h000;
      20'h0339b: out <= 12'h000;
      20'h0339c: out <= 12'h000;
      20'h0339d: out <= 12'h000;
      20'h0339e: out <= 12'h000;
      20'h0339f: out <= 12'h000;
      20'h033a0: out <= 12'h000;
      20'h033a1: out <= 12'h000;
      20'h033a2: out <= 12'h000;
      20'h033a3: out <= 12'h000;
      20'h033a4: out <= 12'h000;
      20'h033a5: out <= 12'h000;
      20'h033a6: out <= 12'h000;
      20'h033a7: out <= 12'h000;
      20'h033a8: out <= 12'h222;
      20'h033a9: out <= 12'h222;
      20'h033aa: out <= 12'h222;
      20'h033ab: out <= 12'h222;
      20'h033ac: out <= 12'h222;
      20'h033ad: out <= 12'h222;
      20'h033ae: out <= 12'h222;
      20'h033af: out <= 12'h222;
      20'h033b0: out <= 12'h222;
      20'h033b1: out <= 12'h222;
      20'h033b2: out <= 12'h222;
      20'h033b3: out <= 12'h222;
      20'h033b4: out <= 12'h222;
      20'h033b5: out <= 12'h222;
      20'h033b6: out <= 12'h222;
      20'h033b7: out <= 12'h222;
      20'h033b8: out <= 12'h000;
      20'h033b9: out <= 12'h000;
      20'h033ba: out <= 12'h000;
      20'h033bb: out <= 12'h000;
      20'h033bc: out <= 12'h000;
      20'h033bd: out <= 12'h000;
      20'h033be: out <= 12'h000;
      20'h033bf: out <= 12'h000;
      20'h033c0: out <= 12'h000;
      20'h033c1: out <= 12'h000;
      20'h033c2: out <= 12'h000;
      20'h033c3: out <= 12'h000;
      20'h033c4: out <= 12'h000;
      20'h033c5: out <= 12'h000;
      20'h033c6: out <= 12'h000;
      20'h033c7: out <= 12'h000;
      20'h033c8: out <= 12'h222;
      20'h033c9: out <= 12'h222;
      20'h033ca: out <= 12'h222;
      20'h033cb: out <= 12'h222;
      20'h033cc: out <= 12'h222;
      20'h033cd: out <= 12'h222;
      20'h033ce: out <= 12'h222;
      20'h033cf: out <= 12'hc7f;
      20'h033d0: out <= 12'hfff;
      20'h033d1: out <= 12'hc7f;
      20'h033d2: out <= 12'h222;
      20'h033d3: out <= 12'h222;
      20'h033d4: out <= 12'h222;
      20'h033d5: out <= 12'h222;
      20'h033d6: out <= 12'h222;
      20'h033d7: out <= 12'h222;
      20'h033d8: out <= 12'h000;
      20'h033d9: out <= 12'h000;
      20'h033da: out <= 12'h000;
      20'h033db: out <= 12'h000;
      20'h033dc: out <= 12'h000;
      20'h033dd: out <= 12'h000;
      20'h033de: out <= 12'h000;
      20'h033df: out <= 12'hc7f;
      20'h033e0: out <= 12'hfff;
      20'h033e1: out <= 12'hc7f;
      20'h033e2: out <= 12'h000;
      20'h033e3: out <= 12'h000;
      20'h033e4: out <= 12'h000;
      20'h033e5: out <= 12'h000;
      20'h033e6: out <= 12'h000;
      20'h033e7: out <= 12'h000;
      20'h033e8: out <= 12'h603;
      20'h033e9: out <= 12'h603;
      20'h033ea: out <= 12'h603;
      20'h033eb: out <= 12'h603;
      20'h033ec: out <= 12'h6af;
      20'h033ed: out <= 12'h4cd;
      20'h033ee: out <= 12'h4cd;
      20'h033ef: out <= 12'h6af;
      20'h033f0: out <= 12'hfff;
      20'h033f1: out <= 12'h4cd;
      20'h033f2: out <= 12'h4cd;
      20'h033f3: out <= 12'hfff;
      20'h033f4: out <= 12'h6af;
      20'h033f5: out <= 12'h4cd;
      20'h033f6: out <= 12'h4cd;
      20'h033f7: out <= 12'h6af;
      20'h033f8: out <= 12'hfff;
      20'h033f9: out <= 12'h4cd;
      20'h033fa: out <= 12'h4cd;
      20'h033fb: out <= 12'hfff;
      20'h033fc: out <= 12'h000;
      20'h033fd: out <= 12'h000;
      20'h033fe: out <= 12'h380;
      20'h033ff: out <= 12'h380;
      20'h03400: out <= 12'h380;
      20'h03401: out <= 12'h380;
      20'h03402: out <= 12'h000;
      20'h03403: out <= 12'h000;
      20'h03404: out <= 12'h000;
      20'h03405: out <= 12'h000;
      20'h03406: out <= 12'h380;
      20'h03407: out <= 12'h380;
      20'h03408: out <= 12'h380;
      20'h03409: out <= 12'h380;
      20'h0340a: out <= 12'h000;
      20'h0340b: out <= 12'h000;
      20'h0340c: out <= 12'h000;
      20'h0340d: out <= 12'h000;
      20'h0340e: out <= 12'hbbb;
      20'h0340f: out <= 12'hfff;
      20'h03410: out <= 12'h000;
      20'h03411: out <= 12'h000;
      20'h03412: out <= 12'hbbb;
      20'h03413: out <= 12'hfff;
      20'h03414: out <= 12'h000;
      20'h03415: out <= 12'h000;
      20'h03416: out <= 12'hbbb;
      20'h03417: out <= 12'hfff;
      20'h03418: out <= 12'h000;
      20'h03419: out <= 12'h000;
      20'h0341a: out <= 12'hbbb;
      20'h0341b: out <= 12'hfff;
      20'h0341c: out <= 12'h000;
      20'h0341d: out <= 12'h000;
      20'h0341e: out <= 12'h000;
      20'h0341f: out <= 12'h000;
      20'h03420: out <= 12'h000;
      20'h03421: out <= 12'h000;
      20'h03422: out <= 12'h000;
      20'h03423: out <= 12'h000;
      20'h03424: out <= 12'h000;
      20'h03425: out <= 12'h000;
      20'h03426: out <= 12'h000;
      20'h03427: out <= 12'h000;
      20'h03428: out <= 12'h000;
      20'h03429: out <= 12'h000;
      20'h0342a: out <= 12'h000;
      20'h0342b: out <= 12'h000;
      20'h0342c: out <= 12'h000;
      20'h0342d: out <= 12'h000;
      20'h0342e: out <= 12'h000;
      20'h0342f: out <= 12'h000;
      20'h03430: out <= 12'h000;
      20'h03431: out <= 12'h000;
      20'h03432: out <= 12'h000;
      20'h03433: out <= 12'h000;
      20'h03434: out <= 12'h000;
      20'h03435: out <= 12'h000;
      20'h03436: out <= 12'h000;
      20'h03437: out <= 12'h000;
      20'h03438: out <= 12'h000;
      20'h03439: out <= 12'h000;
      20'h0343a: out <= 12'h000;
      20'h0343b: out <= 12'h000;
      20'h0343c: out <= 12'h603;
      20'h0343d: out <= 12'h603;
      20'h0343e: out <= 12'h603;
      20'h0343f: out <= 12'h603;
      20'h03440: out <= 12'hb27;
      20'h03441: out <= 12'hb27;
      20'h03442: out <= 12'hb27;
      20'h03443: out <= 12'hb27;
      20'h03444: out <= 12'hb27;
      20'h03445: out <= 12'hb27;
      20'h03446: out <= 12'hb27;
      20'h03447: out <= 12'hb27;
      20'h03448: out <= 12'h000;
      20'h03449: out <= 12'h000;
      20'h0344a: out <= 12'h000;
      20'h0344b: out <= 12'h000;
      20'h0344c: out <= 12'h000;
      20'h0344d: out <= 12'h000;
      20'h0344e: out <= 12'h000;
      20'h0344f: out <= 12'h000;
      20'h03450: out <= 12'h000;
      20'h03451: out <= 12'h000;
      20'h03452: out <= 12'h000;
      20'h03453: out <= 12'h000;
      20'h03454: out <= 12'h000;
      20'h03455: out <= 12'h000;
      20'h03456: out <= 12'h000;
      20'h03457: out <= 12'h000;
      20'h03458: out <= 12'h916;
      20'h03459: out <= 12'h916;
      20'h0345a: out <= 12'h916;
      20'h0345b: out <= 12'h916;
      20'h0345c: out <= 12'h916;
      20'h0345d: out <= 12'h916;
      20'h0345e: out <= 12'h916;
      20'h0345f: out <= 12'h916;
      20'h03460: out <= 12'hd29;
      20'h03461: out <= 12'hd29;
      20'h03462: out <= 12'hd29;
      20'h03463: out <= 12'hd29;
      20'h03464: out <= 12'hd29;
      20'h03465: out <= 12'hd29;
      20'h03466: out <= 12'hd29;
      20'h03467: out <= 12'hd29;
      20'h03468: out <= 12'h000;
      20'h03469: out <= 12'h000;
      20'h0346a: out <= 12'h000;
      20'h0346b: out <= 12'h000;
      20'h0346c: out <= 12'h000;
      20'h0346d: out <= 12'h000;
      20'h0346e: out <= 12'h000;
      20'h0346f: out <= 12'h000;
      20'h03470: out <= 12'h000;
      20'h03471: out <= 12'h000;
      20'h03472: out <= 12'h000;
      20'h03473: out <= 12'h000;
      20'h03474: out <= 12'h000;
      20'h03475: out <= 12'h000;
      20'h03476: out <= 12'h000;
      20'h03477: out <= 12'h000;
      20'h03478: out <= 12'h000;
      20'h03479: out <= 12'h000;
      20'h0347a: out <= 12'h000;
      20'h0347b: out <= 12'h000;
      20'h0347c: out <= 12'h000;
      20'h0347d: out <= 12'h000;
      20'h0347e: out <= 12'h000;
      20'h0347f: out <= 12'h000;
      20'h03480: out <= 12'h000;
      20'h03481: out <= 12'hc7f;
      20'h03482: out <= 12'hfff;
      20'h03483: out <= 12'hc7f;
      20'h03484: out <= 12'hfff;
      20'h03485: out <= 12'hfff;
      20'h03486: out <= 12'hfff;
      20'h03487: out <= 12'hfff;
      20'h03488: out <= 12'hfff;
      20'h03489: out <= 12'hc7f;
      20'h0348a: out <= 12'hc7f;
      20'h0348b: out <= 12'hfff;
      20'h0348c: out <= 12'hc7f;
      20'h0348d: out <= 12'h000;
      20'h0348e: out <= 12'h000;
      20'h0348f: out <= 12'h000;
      20'h03490: out <= 12'h222;
      20'h03491: out <= 12'hc7f;
      20'h03492: out <= 12'hfff;
      20'h03493: out <= 12'hc7f;
      20'h03494: out <= 12'h72f;
      20'h03495: out <= 12'h72f;
      20'h03496: out <= 12'h72f;
      20'h03497: out <= 12'h72f;
      20'h03498: out <= 12'h72f;
      20'h03499: out <= 12'hc7f;
      20'h0349a: out <= 12'hc7f;
      20'h0349b: out <= 12'hfff;
      20'h0349c: out <= 12'hc7f;
      20'h0349d: out <= 12'h222;
      20'h0349e: out <= 12'h222;
      20'h0349f: out <= 12'h222;
      20'h034a0: out <= 12'h000;
      20'h034a1: out <= 12'h000;
      20'h034a2: out <= 12'h000;
      20'h034a3: out <= 12'h000;
      20'h034a4: out <= 12'h000;
      20'h034a5: out <= 12'h000;
      20'h034a6: out <= 12'h000;
      20'h034a7: out <= 12'hc7f;
      20'h034a8: out <= 12'hfff;
      20'h034a9: out <= 12'hc7f;
      20'h034aa: out <= 12'h000;
      20'h034ab: out <= 12'h000;
      20'h034ac: out <= 12'h000;
      20'h034ad: out <= 12'h000;
      20'h034ae: out <= 12'h000;
      20'h034af: out <= 12'h000;
      20'h034b0: out <= 12'h222;
      20'h034b1: out <= 12'h222;
      20'h034b2: out <= 12'h222;
      20'h034b3: out <= 12'h222;
      20'h034b4: out <= 12'h222;
      20'h034b5: out <= 12'h222;
      20'h034b6: out <= 12'h222;
      20'h034b7: out <= 12'hc7f;
      20'h034b8: out <= 12'hfff;
      20'h034b9: out <= 12'hc7f;
      20'h034ba: out <= 12'h222;
      20'h034bb: out <= 12'h222;
      20'h034bc: out <= 12'h222;
      20'h034bd: out <= 12'h222;
      20'h034be: out <= 12'h222;
      20'h034bf: out <= 12'h222;
      20'h034c0: out <= 12'h000;
      20'h034c1: out <= 12'h000;
      20'h034c2: out <= 12'h000;
      20'h034c3: out <= 12'hc7f;
      20'h034c4: out <= 12'hfff;
      20'h034c5: out <= 12'hc7f;
      20'h034c6: out <= 12'hc7f;
      20'h034c7: out <= 12'hfff;
      20'h034c8: out <= 12'hfff;
      20'h034c9: out <= 12'hfff;
      20'h034ca: out <= 12'hfff;
      20'h034cb: out <= 12'hfff;
      20'h034cc: out <= 12'hc7f;
      20'h034cd: out <= 12'hfff;
      20'h034ce: out <= 12'hc7f;
      20'h034cf: out <= 12'h000;
      20'h034d0: out <= 12'h222;
      20'h034d1: out <= 12'h222;
      20'h034d2: out <= 12'h222;
      20'h034d3: out <= 12'hc7f;
      20'h034d4: out <= 12'hfff;
      20'h034d5: out <= 12'hc7f;
      20'h034d6: out <= 12'hc7f;
      20'h034d7: out <= 12'h72f;
      20'h034d8: out <= 12'h72f;
      20'h034d9: out <= 12'h72f;
      20'h034da: out <= 12'h72f;
      20'h034db: out <= 12'h72f;
      20'h034dc: out <= 12'hc7f;
      20'h034dd: out <= 12'hfff;
      20'h034de: out <= 12'hc7f;
      20'h034df: out <= 12'h222;
      20'h034e0: out <= 12'h000;
      20'h034e1: out <= 12'h000;
      20'h034e2: out <= 12'h000;
      20'h034e3: out <= 12'h000;
      20'h034e4: out <= 12'h000;
      20'h034e5: out <= 12'h000;
      20'h034e6: out <= 12'hfff;
      20'h034e7: out <= 12'hfff;
      20'h034e8: out <= 12'hfff;
      20'h034e9: out <= 12'hfff;
      20'h034ea: out <= 12'hfff;
      20'h034eb: out <= 12'h000;
      20'h034ec: out <= 12'h000;
      20'h034ed: out <= 12'h000;
      20'h034ee: out <= 12'h000;
      20'h034ef: out <= 12'h000;
      20'h034f0: out <= 12'h222;
      20'h034f1: out <= 12'h222;
      20'h034f2: out <= 12'h222;
      20'h034f3: out <= 12'h222;
      20'h034f4: out <= 12'h222;
      20'h034f5: out <= 12'h222;
      20'h034f6: out <= 12'h72f;
      20'h034f7: out <= 12'h72f;
      20'h034f8: out <= 12'h72f;
      20'h034f9: out <= 12'h72f;
      20'h034fa: out <= 12'h72f;
      20'h034fb: out <= 12'h222;
      20'h034fc: out <= 12'h222;
      20'h034fd: out <= 12'h222;
      20'h034fe: out <= 12'h222;
      20'h034ff: out <= 12'h222;
      20'h03500: out <= 12'h603;
      20'h03501: out <= 12'h603;
      20'h03502: out <= 12'h603;
      20'h03503: out <= 12'h603;
      20'h03504: out <= 12'h000;
      20'h03505: out <= 12'h000;
      20'h03506: out <= 12'h000;
      20'h03507: out <= 12'h000;
      20'h03508: out <= 12'h000;
      20'h03509: out <= 12'h000;
      20'h0350a: out <= 12'h000;
      20'h0350b: out <= 12'h000;
      20'h0350c: out <= 12'h000;
      20'h0350d: out <= 12'h000;
      20'h0350e: out <= 12'h000;
      20'h0350f: out <= 12'h000;
      20'h03510: out <= 12'h000;
      20'h03511: out <= 12'h000;
      20'h03512: out <= 12'h000;
      20'h03513: out <= 12'h000;
      20'h03514: out <= 12'h000;
      20'h03515: out <= 12'hee9;
      20'h03516: out <= 12'hee9;
      20'h03517: out <= 12'hee9;
      20'h03518: out <= 12'hf87;
      20'h03519: out <= 12'hf87;
      20'h0351a: out <= 12'hf87;
      20'h0351b: out <= 12'hf87;
      20'h0351c: out <= 12'hf87;
      20'h0351d: out <= 12'hf87;
      20'h0351e: out <= 12'hf87;
      20'h0351f: out <= 12'hf87;
      20'h03520: out <= 12'hf87;
      20'h03521: out <= 12'hee9;
      20'h03522: out <= 12'hee9;
      20'h03523: out <= 12'hee9;
      20'h03524: out <= 12'h000;
      20'h03525: out <= 12'h000;
      20'h03526: out <= 12'h000;
      20'h03527: out <= 12'h000;
      20'h03528: out <= 12'h000;
      20'h03529: out <= 12'h000;
      20'h0352a: out <= 12'h000;
      20'h0352b: out <= 12'h000;
      20'h0352c: out <= 12'h000;
      20'h0352d: out <= 12'h000;
      20'h0352e: out <= 12'h000;
      20'h0352f: out <= 12'h000;
      20'h03530: out <= 12'h000;
      20'h03531: out <= 12'h000;
      20'h03532: out <= 12'h000;
      20'h03533: out <= 12'h000;
      20'h03534: out <= 12'h603;
      20'h03535: out <= 12'h603;
      20'h03536: out <= 12'h603;
      20'h03537: out <= 12'h603;
      20'h03538: out <= 12'h603;
      20'h03539: out <= 12'h603;
      20'h0353a: out <= 12'h603;
      20'h0353b: out <= 12'h603;
      20'h0353c: out <= 12'h603;
      20'h0353d: out <= 12'h603;
      20'h0353e: out <= 12'h603;
      20'h0353f: out <= 12'h603;
      20'h03540: out <= 12'h603;
      20'h03541: out <= 12'h603;
      20'h03542: out <= 12'h603;
      20'h03543: out <= 12'h603;
      20'h03544: out <= 12'h603;
      20'h03545: out <= 12'h603;
      20'h03546: out <= 12'h603;
      20'h03547: out <= 12'h603;
      20'h03548: out <= 12'h603;
      20'h03549: out <= 12'h603;
      20'h0354a: out <= 12'h603;
      20'h0354b: out <= 12'h603;
      20'h0354c: out <= 12'h603;
      20'h0354d: out <= 12'h603;
      20'h0354e: out <= 12'h603;
      20'h0354f: out <= 12'h603;
      20'h03550: out <= 12'h603;
      20'h03551: out <= 12'h603;
      20'h03552: out <= 12'h603;
      20'h03553: out <= 12'h603;
      20'h03554: out <= 12'h603;
      20'h03555: out <= 12'h603;
      20'h03556: out <= 12'h603;
      20'h03557: out <= 12'h603;
      20'h03558: out <= 12'hee9;
      20'h03559: out <= 12'hee9;
      20'h0355a: out <= 12'hee9;
      20'h0355b: out <= 12'hee9;
      20'h0355c: out <= 12'hee9;
      20'h0355d: out <= 12'hee9;
      20'h0355e: out <= 12'hee9;
      20'h0355f: out <= 12'hb27;
      20'h03560: out <= 12'hee9;
      20'h03561: out <= 12'hee9;
      20'h03562: out <= 12'hee9;
      20'h03563: out <= 12'hee9;
      20'h03564: out <= 12'hee9;
      20'h03565: out <= 12'hee9;
      20'h03566: out <= 12'hee9;
      20'h03567: out <= 12'hb27;
      20'h03568: out <= 12'hee9;
      20'h03569: out <= 12'hee9;
      20'h0356a: out <= 12'hee9;
      20'h0356b: out <= 12'hee9;
      20'h0356c: out <= 12'hee9;
      20'h0356d: out <= 12'hee9;
      20'h0356e: out <= 12'hee9;
      20'h0356f: out <= 12'hb27;
      20'h03570: out <= 12'hee9;
      20'h03571: out <= 12'hee9;
      20'h03572: out <= 12'hee9;
      20'h03573: out <= 12'hee9;
      20'h03574: out <= 12'hee9;
      20'h03575: out <= 12'hee9;
      20'h03576: out <= 12'hee9;
      20'h03577: out <= 12'hb27;
      20'h03578: out <= 12'hee9;
      20'h03579: out <= 12'hee9;
      20'h0357a: out <= 12'hee9;
      20'h0357b: out <= 12'hee9;
      20'h0357c: out <= 12'hee9;
      20'h0357d: out <= 12'hee9;
      20'h0357e: out <= 12'hee9;
      20'h0357f: out <= 12'hb27;
      20'h03580: out <= 12'hee9;
      20'h03581: out <= 12'hee9;
      20'h03582: out <= 12'hee9;
      20'h03583: out <= 12'hee9;
      20'h03584: out <= 12'hee9;
      20'h03585: out <= 12'hee9;
      20'h03586: out <= 12'hee9;
      20'h03587: out <= 12'hb27;
      20'h03588: out <= 12'hee9;
      20'h03589: out <= 12'hee9;
      20'h0358a: out <= 12'hee9;
      20'h0358b: out <= 12'hee9;
      20'h0358c: out <= 12'hee9;
      20'h0358d: out <= 12'hee9;
      20'h0358e: out <= 12'hee9;
      20'h0358f: out <= 12'hb27;
      20'h03590: out <= 12'hee9;
      20'h03591: out <= 12'hee9;
      20'h03592: out <= 12'hee9;
      20'h03593: out <= 12'hee9;
      20'h03594: out <= 12'hee9;
      20'h03595: out <= 12'hee9;
      20'h03596: out <= 12'hee9;
      20'h03597: out <= 12'hb27;
      20'h03598: out <= 12'h000;
      20'h03599: out <= 12'h72f;
      20'h0359a: out <= 12'hfff;
      20'h0359b: out <= 12'hfff;
      20'h0359c: out <= 12'hc7f;
      20'h0359d: out <= 12'hc7f;
      20'h0359e: out <= 12'hc7f;
      20'h0359f: out <= 12'hc7f;
      20'h035a0: out <= 12'hc7f;
      20'h035a1: out <= 12'hfff;
      20'h035a2: out <= 12'h72f;
      20'h035a3: out <= 12'hfff;
      20'h035a4: out <= 12'h72f;
      20'h035a5: out <= 12'h000;
      20'h035a6: out <= 12'h000;
      20'h035a7: out <= 12'h000;
      20'h035a8: out <= 12'h222;
      20'h035a9: out <= 12'h72f;
      20'h035aa: out <= 12'hfff;
      20'h035ab: out <= 12'h72f;
      20'h035ac: out <= 12'hc7f;
      20'h035ad: out <= 12'hc7f;
      20'h035ae: out <= 12'hc7f;
      20'h035af: out <= 12'hc7f;
      20'h035b0: out <= 12'hc7f;
      20'h035b1: out <= 12'h72f;
      20'h035b2: out <= 12'h72f;
      20'h035b3: out <= 12'hfff;
      20'h035b4: out <= 12'h72f;
      20'h035b5: out <= 12'h222;
      20'h035b6: out <= 12'h222;
      20'h035b7: out <= 12'h222;
      20'h035b8: out <= 12'h000;
      20'h035b9: out <= 12'h000;
      20'h035ba: out <= 12'h000;
      20'h035bb: out <= 12'h000;
      20'h035bc: out <= 12'h000;
      20'h035bd: out <= 12'h000;
      20'h035be: out <= 12'h000;
      20'h035bf: out <= 12'h72f;
      20'h035c0: out <= 12'hfff;
      20'h035c1: out <= 12'h72f;
      20'h035c2: out <= 12'h000;
      20'h035c3: out <= 12'h000;
      20'h035c4: out <= 12'h000;
      20'h035c5: out <= 12'h000;
      20'h035c6: out <= 12'h000;
      20'h035c7: out <= 12'h000;
      20'h035c8: out <= 12'h222;
      20'h035c9: out <= 12'h222;
      20'h035ca: out <= 12'h222;
      20'h035cb: out <= 12'h222;
      20'h035cc: out <= 12'h222;
      20'h035cd: out <= 12'h222;
      20'h035ce: out <= 12'h222;
      20'h035cf: out <= 12'h72f;
      20'h035d0: out <= 12'hfff;
      20'h035d1: out <= 12'h72f;
      20'h035d2: out <= 12'h222;
      20'h035d3: out <= 12'h222;
      20'h035d4: out <= 12'h222;
      20'h035d5: out <= 12'h222;
      20'h035d6: out <= 12'h222;
      20'h035d7: out <= 12'h222;
      20'h035d8: out <= 12'h000;
      20'h035d9: out <= 12'h000;
      20'h035da: out <= 12'h000;
      20'h035db: out <= 12'h72f;
      20'h035dc: out <= 12'hfff;
      20'h035dd: out <= 12'h72f;
      20'h035de: out <= 12'hfff;
      20'h035df: out <= 12'hc7f;
      20'h035e0: out <= 12'hc7f;
      20'h035e1: out <= 12'hc7f;
      20'h035e2: out <= 12'hc7f;
      20'h035e3: out <= 12'hc7f;
      20'h035e4: out <= 12'hfff;
      20'h035e5: out <= 12'hfff;
      20'h035e6: out <= 12'h72f;
      20'h035e7: out <= 12'h000;
      20'h035e8: out <= 12'h222;
      20'h035e9: out <= 12'h222;
      20'h035ea: out <= 12'h222;
      20'h035eb: out <= 12'h72f;
      20'h035ec: out <= 12'hfff;
      20'h035ed: out <= 12'h72f;
      20'h035ee: out <= 12'h72f;
      20'h035ef: out <= 12'hc7f;
      20'h035f0: out <= 12'hc7f;
      20'h035f1: out <= 12'hc7f;
      20'h035f2: out <= 12'hc7f;
      20'h035f3: out <= 12'hc7f;
      20'h035f4: out <= 12'h72f;
      20'h035f5: out <= 12'hfff;
      20'h035f6: out <= 12'h72f;
      20'h035f7: out <= 12'h222;
      20'h035f8: out <= 12'h000;
      20'h035f9: out <= 12'hc7f;
      20'h035fa: out <= 12'h72f;
      20'h035fb: out <= 12'hc7f;
      20'h035fc: out <= 12'hfff;
      20'h035fd: out <= 12'hfff;
      20'h035fe: out <= 12'hc7f;
      20'h035ff: out <= 12'hc7f;
      20'h03600: out <= 12'hc7f;
      20'h03601: out <= 12'hc7f;
      20'h03602: out <= 12'hc7f;
      20'h03603: out <= 12'hfff;
      20'h03604: out <= 12'hfff;
      20'h03605: out <= 12'hc7f;
      20'h03606: out <= 12'h72f;
      20'h03607: out <= 12'hc7f;
      20'h03608: out <= 12'h222;
      20'h03609: out <= 12'hc7f;
      20'h0360a: out <= 12'h72f;
      20'h0360b: out <= 12'hc7f;
      20'h0360c: out <= 12'h72f;
      20'h0360d: out <= 12'h72f;
      20'h0360e: out <= 12'hc7f;
      20'h0360f: out <= 12'hc7f;
      20'h03610: out <= 12'hc7f;
      20'h03611: out <= 12'hc7f;
      20'h03612: out <= 12'hc7f;
      20'h03613: out <= 12'h72f;
      20'h03614: out <= 12'h72f;
      20'h03615: out <= 12'hc7f;
      20'h03616: out <= 12'h72f;
      20'h03617: out <= 12'hc7f;
      20'h03618: out <= 12'h603;
      20'h03619: out <= 12'h603;
      20'h0361a: out <= 12'h603;
      20'h0361b: out <= 12'h603;
      20'h0361c: out <= 12'h000;
      20'h0361d: out <= 12'h000;
      20'h0361e: out <= 12'hee9;
      20'h0361f: out <= 12'hb27;
      20'h03620: out <= 12'hb27;
      20'h03621: out <= 12'hb27;
      20'h03622: out <= 12'hb27;
      20'h03623: out <= 12'hb27;
      20'h03624: out <= 12'hb27;
      20'h03625: out <= 12'hb27;
      20'h03626: out <= 12'hb27;
      20'h03627: out <= 12'hb27;
      20'h03628: out <= 12'hb27;
      20'h03629: out <= 12'hb27;
      20'h0362a: out <= 12'hee9;
      20'h0362b: out <= 12'h000;
      20'h0362c: out <= 12'h000;
      20'h0362d: out <= 12'hee9;
      20'h0362e: out <= 12'hf87;
      20'h0362f: out <= 12'hf87;
      20'h03630: out <= 12'hee9;
      20'h03631: out <= 12'hb27;
      20'h03632: out <= 12'hb27;
      20'h03633: out <= 12'hb27;
      20'h03634: out <= 12'hb27;
      20'h03635: out <= 12'hb27;
      20'h03636: out <= 12'hb27;
      20'h03637: out <= 12'hb27;
      20'h03638: out <= 12'hee9;
      20'h03639: out <= 12'hf87;
      20'h0363a: out <= 12'hf87;
      20'h0363b: out <= 12'hb27;
      20'h0363c: out <= 12'h000;
      20'h0363d: out <= 12'h000;
      20'h0363e: out <= 12'h000;
      20'h0363f: out <= 12'h000;
      20'h03640: out <= 12'hee9;
      20'h03641: out <= 12'h000;
      20'h03642: out <= 12'h000;
      20'h03643: out <= 12'h000;
      20'h03644: out <= 12'h000;
      20'h03645: out <= 12'h000;
      20'h03646: out <= 12'h000;
      20'h03647: out <= 12'h000;
      20'h03648: out <= 12'h000;
      20'h03649: out <= 12'h000;
      20'h0364a: out <= 12'h000;
      20'h0364b: out <= 12'h000;
      20'h0364c: out <= 12'h603;
      20'h0364d: out <= 12'h603;
      20'h0364e: out <= 12'h603;
      20'h0364f: out <= 12'h603;
      20'h03650: out <= 12'h603;
      20'h03651: out <= 12'h603;
      20'h03652: out <= 12'h603;
      20'h03653: out <= 12'h603;
      20'h03654: out <= 12'h603;
      20'h03655: out <= 12'h603;
      20'h03656: out <= 12'h603;
      20'h03657: out <= 12'h603;
      20'h03658: out <= 12'h603;
      20'h03659: out <= 12'h603;
      20'h0365a: out <= 12'h603;
      20'h0365b: out <= 12'h603;
      20'h0365c: out <= 12'h603;
      20'h0365d: out <= 12'h603;
      20'h0365e: out <= 12'h603;
      20'h0365f: out <= 12'h603;
      20'h03660: out <= 12'h603;
      20'h03661: out <= 12'h603;
      20'h03662: out <= 12'h603;
      20'h03663: out <= 12'h603;
      20'h03664: out <= 12'h603;
      20'h03665: out <= 12'h603;
      20'h03666: out <= 12'h603;
      20'h03667: out <= 12'h603;
      20'h03668: out <= 12'h603;
      20'h03669: out <= 12'h603;
      20'h0366a: out <= 12'h603;
      20'h0366b: out <= 12'h603;
      20'h0366c: out <= 12'h603;
      20'h0366d: out <= 12'h603;
      20'h0366e: out <= 12'h603;
      20'h0366f: out <= 12'h603;
      20'h03670: out <= 12'hee9;
      20'h03671: out <= 12'hf87;
      20'h03672: out <= 12'hf87;
      20'h03673: out <= 12'hf87;
      20'h03674: out <= 12'hf87;
      20'h03675: out <= 12'hf87;
      20'h03676: out <= 12'hf87;
      20'h03677: out <= 12'hb27;
      20'h03678: out <= 12'hee9;
      20'h03679: out <= 12'hf87;
      20'h0367a: out <= 12'hf87;
      20'h0367b: out <= 12'hf87;
      20'h0367c: out <= 12'hf87;
      20'h0367d: out <= 12'hf87;
      20'h0367e: out <= 12'hf87;
      20'h0367f: out <= 12'hb27;
      20'h03680: out <= 12'hee9;
      20'h03681: out <= 12'hf87;
      20'h03682: out <= 12'hf87;
      20'h03683: out <= 12'hf87;
      20'h03684: out <= 12'hf87;
      20'h03685: out <= 12'hf87;
      20'h03686: out <= 12'hf87;
      20'h03687: out <= 12'hb27;
      20'h03688: out <= 12'hee9;
      20'h03689: out <= 12'hf87;
      20'h0368a: out <= 12'hf87;
      20'h0368b: out <= 12'hf87;
      20'h0368c: out <= 12'hf87;
      20'h0368d: out <= 12'hf87;
      20'h0368e: out <= 12'hf87;
      20'h0368f: out <= 12'hb27;
      20'h03690: out <= 12'hee9;
      20'h03691: out <= 12'hf87;
      20'h03692: out <= 12'hf87;
      20'h03693: out <= 12'hf87;
      20'h03694: out <= 12'hf87;
      20'h03695: out <= 12'hf87;
      20'h03696: out <= 12'hf87;
      20'h03697: out <= 12'hb27;
      20'h03698: out <= 12'hee9;
      20'h03699: out <= 12'hf87;
      20'h0369a: out <= 12'hf87;
      20'h0369b: out <= 12'hf87;
      20'h0369c: out <= 12'hf87;
      20'h0369d: out <= 12'hf87;
      20'h0369e: out <= 12'hf87;
      20'h0369f: out <= 12'hb27;
      20'h036a0: out <= 12'hee9;
      20'h036a1: out <= 12'hf87;
      20'h036a2: out <= 12'hf87;
      20'h036a3: out <= 12'hf87;
      20'h036a4: out <= 12'hf87;
      20'h036a5: out <= 12'hf87;
      20'h036a6: out <= 12'hf87;
      20'h036a7: out <= 12'hb27;
      20'h036a8: out <= 12'hee9;
      20'h036a9: out <= 12'hf87;
      20'h036aa: out <= 12'hf87;
      20'h036ab: out <= 12'hf87;
      20'h036ac: out <= 12'hf87;
      20'h036ad: out <= 12'hf87;
      20'h036ae: out <= 12'hf87;
      20'h036af: out <= 12'hb27;
      20'h036b0: out <= 12'h000;
      20'h036b1: out <= 12'hc7f;
      20'h036b2: out <= 12'hfff;
      20'h036b3: out <= 12'hc7f;
      20'h036b4: out <= 12'h72f;
      20'h036b5: out <= 12'h72f;
      20'h036b6: out <= 12'h72f;
      20'h036b7: out <= 12'h72f;
      20'h036b8: out <= 12'h72f;
      20'h036b9: out <= 12'hc7f;
      20'h036ba: out <= 12'hfff;
      20'h036bb: out <= 12'hfff;
      20'h036bc: out <= 12'hc7f;
      20'h036bd: out <= 12'h000;
      20'h036be: out <= 12'h000;
      20'h036bf: out <= 12'h000;
      20'h036c0: out <= 12'h222;
      20'h036c1: out <= 12'hc7f;
      20'h036c2: out <= 12'hfff;
      20'h036c3: out <= 12'hc7f;
      20'h036c4: out <= 12'hfff;
      20'h036c5: out <= 12'hfff;
      20'h036c6: out <= 12'hfff;
      20'h036c7: out <= 12'hfff;
      20'h036c8: out <= 12'hfff;
      20'h036c9: out <= 12'hc7f;
      20'h036ca: out <= 12'h72f;
      20'h036cb: out <= 12'hfff;
      20'h036cc: out <= 12'hc7f;
      20'h036cd: out <= 12'h222;
      20'h036ce: out <= 12'h222;
      20'h036cf: out <= 12'h222;
      20'h036d0: out <= 12'h000;
      20'h036d1: out <= 12'h000;
      20'h036d2: out <= 12'h000;
      20'h036d3: out <= 12'h000;
      20'h036d4: out <= 12'h000;
      20'h036d5: out <= 12'h000;
      20'h036d6: out <= 12'h000;
      20'h036d7: out <= 12'h72f;
      20'h036d8: out <= 12'hfff;
      20'h036d9: out <= 12'h72f;
      20'h036da: out <= 12'h000;
      20'h036db: out <= 12'h000;
      20'h036dc: out <= 12'h000;
      20'h036dd: out <= 12'h000;
      20'h036de: out <= 12'h000;
      20'h036df: out <= 12'h000;
      20'h036e0: out <= 12'h222;
      20'h036e1: out <= 12'h222;
      20'h036e2: out <= 12'h222;
      20'h036e3: out <= 12'h222;
      20'h036e4: out <= 12'h222;
      20'h036e5: out <= 12'h222;
      20'h036e6: out <= 12'h222;
      20'h036e7: out <= 12'h72f;
      20'h036e8: out <= 12'hfff;
      20'h036e9: out <= 12'h72f;
      20'h036ea: out <= 12'h222;
      20'h036eb: out <= 12'h222;
      20'h036ec: out <= 12'h222;
      20'h036ed: out <= 12'h222;
      20'h036ee: out <= 12'h222;
      20'h036ef: out <= 12'h222;
      20'h036f0: out <= 12'h000;
      20'h036f1: out <= 12'h000;
      20'h036f2: out <= 12'h000;
      20'h036f3: out <= 12'hc7f;
      20'h036f4: out <= 12'hfff;
      20'h036f5: out <= 12'hfff;
      20'h036f6: out <= 12'hc7f;
      20'h036f7: out <= 12'h72f;
      20'h036f8: out <= 12'h72f;
      20'h036f9: out <= 12'h72f;
      20'h036fa: out <= 12'h72f;
      20'h036fb: out <= 12'h72f;
      20'h036fc: out <= 12'hc7f;
      20'h036fd: out <= 12'hfff;
      20'h036fe: out <= 12'hc7f;
      20'h036ff: out <= 12'h000;
      20'h03700: out <= 12'h222;
      20'h03701: out <= 12'h222;
      20'h03702: out <= 12'h222;
      20'h03703: out <= 12'hc7f;
      20'h03704: out <= 12'hfff;
      20'h03705: out <= 12'h72f;
      20'h03706: out <= 12'hc7f;
      20'h03707: out <= 12'hfff;
      20'h03708: out <= 12'hfff;
      20'h03709: out <= 12'hfff;
      20'h0370a: out <= 12'hfff;
      20'h0370b: out <= 12'hfff;
      20'h0370c: out <= 12'hc7f;
      20'h0370d: out <= 12'hfff;
      20'h0370e: out <= 12'hc7f;
      20'h0370f: out <= 12'h222;
      20'h03710: out <= 12'h000;
      20'h03711: out <= 12'hfff;
      20'h03712: out <= 12'hfff;
      20'h03713: out <= 12'hfff;
      20'h03714: out <= 12'hc7f;
      20'h03715: out <= 12'hc7f;
      20'h03716: out <= 12'h72f;
      20'h03717: out <= 12'h72f;
      20'h03718: out <= 12'h72f;
      20'h03719: out <= 12'h72f;
      20'h0371a: out <= 12'h72f;
      20'h0371b: out <= 12'hc7f;
      20'h0371c: out <= 12'hc7f;
      20'h0371d: out <= 12'hfff;
      20'h0371e: out <= 12'hfff;
      20'h0371f: out <= 12'hfff;
      20'h03720: out <= 12'h222;
      20'h03721: out <= 12'hfff;
      20'h03722: out <= 12'hfff;
      20'h03723: out <= 12'hfff;
      20'h03724: out <= 12'hc7f;
      20'h03725: out <= 12'hc7f;
      20'h03726: out <= 12'hfff;
      20'h03727: out <= 12'hfff;
      20'h03728: out <= 12'hfff;
      20'h03729: out <= 12'hfff;
      20'h0372a: out <= 12'hfff;
      20'h0372b: out <= 12'hc7f;
      20'h0372c: out <= 12'hc7f;
      20'h0372d: out <= 12'hfff;
      20'h0372e: out <= 12'hfff;
      20'h0372f: out <= 12'hfff;
      20'h03730: out <= 12'h603;
      20'h03731: out <= 12'h603;
      20'h03732: out <= 12'h603;
      20'h03733: out <= 12'h603;
      20'h03734: out <= 12'h000;
      20'h03735: out <= 12'h000;
      20'h03736: out <= 12'hb27;
      20'h03737: out <= 12'hb27;
      20'h03738: out <= 12'hf87;
      20'h03739: out <= 12'hf87;
      20'h0373a: out <= 12'hf87;
      20'h0373b: out <= 12'hf87;
      20'h0373c: out <= 12'hf87;
      20'h0373d: out <= 12'hf87;
      20'h0373e: out <= 12'hf87;
      20'h0373f: out <= 12'hf87;
      20'h03740: out <= 12'hf87;
      20'h03741: out <= 12'hb27;
      20'h03742: out <= 12'hb27;
      20'h03743: out <= 12'h000;
      20'h03744: out <= 12'h000;
      20'h03745: out <= 12'hee9;
      20'h03746: out <= 12'hf87;
      20'h03747: out <= 12'hb27;
      20'h03748: out <= 12'hf87;
      20'h03749: out <= 12'hee9;
      20'h0374a: out <= 12'hf87;
      20'h0374b: out <= 12'hf87;
      20'h0374c: out <= 12'hf87;
      20'h0374d: out <= 12'hf87;
      20'h0374e: out <= 12'hf87;
      20'h0374f: out <= 12'hee9;
      20'h03750: out <= 12'hf87;
      20'h03751: out <= 12'hb27;
      20'h03752: out <= 12'hf87;
      20'h03753: out <= 12'hb27;
      20'h03754: out <= 12'h000;
      20'h03755: out <= 12'h000;
      20'h03756: out <= 12'h000;
      20'h03757: out <= 12'h000;
      20'h03758: out <= 12'h000;
      20'h03759: out <= 12'hee9;
      20'h0375a: out <= 12'hf87;
      20'h0375b: out <= 12'h000;
      20'h0375c: out <= 12'h000;
      20'h0375d: out <= 12'h000;
      20'h0375e: out <= 12'h000;
      20'h0375f: out <= 12'h000;
      20'h03760: out <= 12'h000;
      20'h03761: out <= 12'h000;
      20'h03762: out <= 12'h000;
      20'h03763: out <= 12'h000;
      20'h03764: out <= 12'h603;
      20'h03765: out <= 12'h603;
      20'h03766: out <= 12'h603;
      20'h03767: out <= 12'h603;
      20'h03768: out <= 12'h603;
      20'h03769: out <= 12'h603;
      20'h0376a: out <= 12'h603;
      20'h0376b: out <= 12'h603;
      20'h0376c: out <= 12'h603;
      20'h0376d: out <= 12'h603;
      20'h0376e: out <= 12'h603;
      20'h0376f: out <= 12'h603;
      20'h03770: out <= 12'h603;
      20'h03771: out <= 12'h603;
      20'h03772: out <= 12'h603;
      20'h03773: out <= 12'h603;
      20'h03774: out <= 12'h603;
      20'h03775: out <= 12'h603;
      20'h03776: out <= 12'h603;
      20'h03777: out <= 12'h603;
      20'h03778: out <= 12'h603;
      20'h03779: out <= 12'h603;
      20'h0377a: out <= 12'h603;
      20'h0377b: out <= 12'h603;
      20'h0377c: out <= 12'h603;
      20'h0377d: out <= 12'h603;
      20'h0377e: out <= 12'h603;
      20'h0377f: out <= 12'h603;
      20'h03780: out <= 12'h603;
      20'h03781: out <= 12'h603;
      20'h03782: out <= 12'h603;
      20'h03783: out <= 12'h603;
      20'h03784: out <= 12'h603;
      20'h03785: out <= 12'h603;
      20'h03786: out <= 12'h603;
      20'h03787: out <= 12'h603;
      20'h03788: out <= 12'hee9;
      20'h03789: out <= 12'hf87;
      20'h0378a: out <= 12'hee9;
      20'h0378b: out <= 12'hee9;
      20'h0378c: out <= 12'hee9;
      20'h0378d: out <= 12'hb27;
      20'h0378e: out <= 12'hf87;
      20'h0378f: out <= 12'hb27;
      20'h03790: out <= 12'hee9;
      20'h03791: out <= 12'hf87;
      20'h03792: out <= 12'hee9;
      20'h03793: out <= 12'hee9;
      20'h03794: out <= 12'hee9;
      20'h03795: out <= 12'hb27;
      20'h03796: out <= 12'hf87;
      20'h03797: out <= 12'hb27;
      20'h03798: out <= 12'hee9;
      20'h03799: out <= 12'hf87;
      20'h0379a: out <= 12'hee9;
      20'h0379b: out <= 12'hee9;
      20'h0379c: out <= 12'hee9;
      20'h0379d: out <= 12'hb27;
      20'h0379e: out <= 12'hf87;
      20'h0379f: out <= 12'hb27;
      20'h037a0: out <= 12'hee9;
      20'h037a1: out <= 12'hf87;
      20'h037a2: out <= 12'hee9;
      20'h037a3: out <= 12'hee9;
      20'h037a4: out <= 12'hee9;
      20'h037a5: out <= 12'hb27;
      20'h037a6: out <= 12'hf87;
      20'h037a7: out <= 12'hb27;
      20'h037a8: out <= 12'hee9;
      20'h037a9: out <= 12'hf87;
      20'h037aa: out <= 12'hee9;
      20'h037ab: out <= 12'hee9;
      20'h037ac: out <= 12'hee9;
      20'h037ad: out <= 12'hb27;
      20'h037ae: out <= 12'hf87;
      20'h037af: out <= 12'hb27;
      20'h037b0: out <= 12'hee9;
      20'h037b1: out <= 12'hf87;
      20'h037b2: out <= 12'hee9;
      20'h037b3: out <= 12'hee9;
      20'h037b4: out <= 12'hee9;
      20'h037b5: out <= 12'hb27;
      20'h037b6: out <= 12'hf87;
      20'h037b7: out <= 12'hb27;
      20'h037b8: out <= 12'hee9;
      20'h037b9: out <= 12'hf87;
      20'h037ba: out <= 12'hee9;
      20'h037bb: out <= 12'hee9;
      20'h037bc: out <= 12'hee9;
      20'h037bd: out <= 12'hb27;
      20'h037be: out <= 12'hf87;
      20'h037bf: out <= 12'hb27;
      20'h037c0: out <= 12'hee9;
      20'h037c1: out <= 12'hf87;
      20'h037c2: out <= 12'hee9;
      20'h037c3: out <= 12'hee9;
      20'h037c4: out <= 12'hee9;
      20'h037c5: out <= 12'hb27;
      20'h037c6: out <= 12'hf87;
      20'h037c7: out <= 12'hb27;
      20'h037c8: out <= 12'h000;
      20'h037c9: out <= 12'hfff;
      20'h037ca: out <= 12'hc7f;
      20'h037cb: out <= 12'h72f;
      20'h037cc: out <= 12'h72f;
      20'h037cd: out <= 12'h72f;
      20'h037ce: out <= 12'h72f;
      20'h037cf: out <= 12'h72f;
      20'h037d0: out <= 12'h72f;
      20'h037d1: out <= 12'h72f;
      20'h037d2: out <= 12'hc7f;
      20'h037d3: out <= 12'hfff;
      20'h037d4: out <= 12'h000;
      20'h037d5: out <= 12'h000;
      20'h037d6: out <= 12'h000;
      20'h037d7: out <= 12'h000;
      20'h037d8: out <= 12'h222;
      20'h037d9: out <= 12'h72f;
      20'h037da: out <= 12'hc7f;
      20'h037db: out <= 12'hfff;
      20'h037dc: out <= 12'h72f;
      20'h037dd: out <= 12'h72f;
      20'h037de: out <= 12'h72f;
      20'h037df: out <= 12'h72f;
      20'h037e0: out <= 12'h72f;
      20'h037e1: out <= 12'hfff;
      20'h037e2: out <= 12'hc7f;
      20'h037e3: out <= 12'h72f;
      20'h037e4: out <= 12'h222;
      20'h037e5: out <= 12'h222;
      20'h037e6: out <= 12'h222;
      20'h037e7: out <= 12'h222;
      20'h037e8: out <= 12'h000;
      20'h037e9: out <= 12'hc7f;
      20'h037ea: out <= 12'h72f;
      20'h037eb: out <= 12'hc7f;
      20'h037ec: out <= 12'h000;
      20'h037ed: out <= 12'h000;
      20'h037ee: out <= 12'hfff;
      20'h037ef: out <= 12'hfff;
      20'h037f0: out <= 12'hfff;
      20'h037f1: out <= 12'hfff;
      20'h037f2: out <= 12'hfff;
      20'h037f3: out <= 12'h000;
      20'h037f4: out <= 12'h000;
      20'h037f5: out <= 12'hc7f;
      20'h037f6: out <= 12'h72f;
      20'h037f7: out <= 12'hc7f;
      20'h037f8: out <= 12'h222;
      20'h037f9: out <= 12'hc7f;
      20'h037fa: out <= 12'h72f;
      20'h037fb: out <= 12'hc7f;
      20'h037fc: out <= 12'h222;
      20'h037fd: out <= 12'h222;
      20'h037fe: out <= 12'h72f;
      20'h037ff: out <= 12'h72f;
      20'h03800: out <= 12'h72f;
      20'h03801: out <= 12'h72f;
      20'h03802: out <= 12'h72f;
      20'h03803: out <= 12'h222;
      20'h03804: out <= 12'h222;
      20'h03805: out <= 12'hc7f;
      20'h03806: out <= 12'h72f;
      20'h03807: out <= 12'hc7f;
      20'h03808: out <= 12'h000;
      20'h03809: out <= 12'h000;
      20'h0380a: out <= 12'h000;
      20'h0380b: out <= 12'h000;
      20'h0380c: out <= 12'hfff;
      20'h0380d: out <= 12'hc7f;
      20'h0380e: out <= 12'h72f;
      20'h0380f: out <= 12'h72f;
      20'h03810: out <= 12'h72f;
      20'h03811: out <= 12'h72f;
      20'h03812: out <= 12'h72f;
      20'h03813: out <= 12'h72f;
      20'h03814: out <= 12'h72f;
      20'h03815: out <= 12'hc7f;
      20'h03816: out <= 12'hfff;
      20'h03817: out <= 12'h000;
      20'h03818: out <= 12'h222;
      20'h03819: out <= 12'h222;
      20'h0381a: out <= 12'h222;
      20'h0381b: out <= 12'h222;
      20'h0381c: out <= 12'h72f;
      20'h0381d: out <= 12'hc7f;
      20'h0381e: out <= 12'hfff;
      20'h0381f: out <= 12'h72f;
      20'h03820: out <= 12'h72f;
      20'h03821: out <= 12'h72f;
      20'h03822: out <= 12'h72f;
      20'h03823: out <= 12'h72f;
      20'h03824: out <= 12'hfff;
      20'h03825: out <= 12'hc7f;
      20'h03826: out <= 12'h72f;
      20'h03827: out <= 12'h222;
      20'h03828: out <= 12'h000;
      20'h03829: out <= 12'hc7f;
      20'h0382a: out <= 12'hfff;
      20'h0382b: out <= 12'hc7f;
      20'h0382c: out <= 12'h72f;
      20'h0382d: out <= 12'h72f;
      20'h0382e: out <= 12'hc7f;
      20'h0382f: out <= 12'hfff;
      20'h03830: out <= 12'hfff;
      20'h03831: out <= 12'hfff;
      20'h03832: out <= 12'hc7f;
      20'h03833: out <= 12'h72f;
      20'h03834: out <= 12'h72f;
      20'h03835: out <= 12'hc7f;
      20'h03836: out <= 12'hfff;
      20'h03837: out <= 12'hc7f;
      20'h03838: out <= 12'h222;
      20'h03839: out <= 12'hc7f;
      20'h0383a: out <= 12'h72f;
      20'h0383b: out <= 12'hc7f;
      20'h0383c: out <= 12'hfff;
      20'h0383d: out <= 12'hfff;
      20'h0383e: out <= 12'hc7f;
      20'h0383f: out <= 12'hfff;
      20'h03840: out <= 12'hfff;
      20'h03841: out <= 12'hfff;
      20'h03842: out <= 12'hc7f;
      20'h03843: out <= 12'hfff;
      20'h03844: out <= 12'hfff;
      20'h03845: out <= 12'hc7f;
      20'h03846: out <= 12'h72f;
      20'h03847: out <= 12'hc7f;
      20'h03848: out <= 12'h603;
      20'h03849: out <= 12'h603;
      20'h0384a: out <= 12'h603;
      20'h0384b: out <= 12'h603;
      20'h0384c: out <= 12'h000;
      20'h0384d: out <= 12'h000;
      20'h0384e: out <= 12'hb27;
      20'h0384f: out <= 12'hf87;
      20'h03850: out <= 12'hf87;
      20'h03851: out <= 12'hee9;
      20'h03852: out <= 12'hee9;
      20'h03853: out <= 12'hee9;
      20'h03854: out <= 12'hee9;
      20'h03855: out <= 12'hee9;
      20'h03856: out <= 12'hee9;
      20'h03857: out <= 12'hee9;
      20'h03858: out <= 12'hf87;
      20'h03859: out <= 12'hf87;
      20'h0385a: out <= 12'hb27;
      20'h0385b: out <= 12'h000;
      20'h0385c: out <= 12'h000;
      20'h0385d: out <= 12'hf87;
      20'h0385e: out <= 12'hb27;
      20'h0385f: out <= 12'hf87;
      20'h03860: out <= 12'hf87;
      20'h03861: out <= 12'hf87;
      20'h03862: out <= 12'hee9;
      20'h03863: out <= 12'hf87;
      20'h03864: out <= 12'hf87;
      20'h03865: out <= 12'hf87;
      20'h03866: out <= 12'hee9;
      20'h03867: out <= 12'hf87;
      20'h03868: out <= 12'hf87;
      20'h03869: out <= 12'hf87;
      20'h0386a: out <= 12'hb27;
      20'h0386b: out <= 12'hf87;
      20'h0386c: out <= 12'h000;
      20'h0386d: out <= 12'h000;
      20'h0386e: out <= 12'h000;
      20'h0386f: out <= 12'hf87;
      20'h03870: out <= 12'hf87;
      20'h03871: out <= 12'hf87;
      20'h03872: out <= 12'hee9;
      20'h03873: out <= 12'h000;
      20'h03874: out <= 12'h000;
      20'h03875: out <= 12'h000;
      20'h03876: out <= 12'hee9;
      20'h03877: out <= 12'hf87;
      20'h03878: out <= 12'h000;
      20'h03879: out <= 12'h000;
      20'h0387a: out <= 12'h000;
      20'h0387b: out <= 12'h000;
      20'h0387c: out <= 12'h603;
      20'h0387d: out <= 12'h603;
      20'h0387e: out <= 12'h603;
      20'h0387f: out <= 12'h603;
      20'h03880: out <= 12'h603;
      20'h03881: out <= 12'h603;
      20'h03882: out <= 12'h603;
      20'h03883: out <= 12'h603;
      20'h03884: out <= 12'h603;
      20'h03885: out <= 12'h603;
      20'h03886: out <= 12'h603;
      20'h03887: out <= 12'h603;
      20'h03888: out <= 12'h603;
      20'h03889: out <= 12'h603;
      20'h0388a: out <= 12'h603;
      20'h0388b: out <= 12'h603;
      20'h0388c: out <= 12'h603;
      20'h0388d: out <= 12'h603;
      20'h0388e: out <= 12'h603;
      20'h0388f: out <= 12'h603;
      20'h03890: out <= 12'h603;
      20'h03891: out <= 12'h603;
      20'h03892: out <= 12'h603;
      20'h03893: out <= 12'h603;
      20'h03894: out <= 12'h603;
      20'h03895: out <= 12'h603;
      20'h03896: out <= 12'h603;
      20'h03897: out <= 12'h603;
      20'h03898: out <= 12'h603;
      20'h03899: out <= 12'h603;
      20'h0389a: out <= 12'h603;
      20'h0389b: out <= 12'h603;
      20'h0389c: out <= 12'h603;
      20'h0389d: out <= 12'h603;
      20'h0389e: out <= 12'h603;
      20'h0389f: out <= 12'h603;
      20'h038a0: out <= 12'hee9;
      20'h038a1: out <= 12'hf87;
      20'h038a2: out <= 12'hee9;
      20'h038a3: out <= 12'hf87;
      20'h038a4: out <= 12'hf87;
      20'h038a5: out <= 12'hb27;
      20'h038a6: out <= 12'hf87;
      20'h038a7: out <= 12'hb27;
      20'h038a8: out <= 12'hee9;
      20'h038a9: out <= 12'hf87;
      20'h038aa: out <= 12'hee9;
      20'h038ab: out <= 12'hf87;
      20'h038ac: out <= 12'hf87;
      20'h038ad: out <= 12'hb27;
      20'h038ae: out <= 12'hf87;
      20'h038af: out <= 12'hb27;
      20'h038b0: out <= 12'hee9;
      20'h038b1: out <= 12'hf87;
      20'h038b2: out <= 12'hee9;
      20'h038b3: out <= 12'hf87;
      20'h038b4: out <= 12'hf87;
      20'h038b5: out <= 12'hb27;
      20'h038b6: out <= 12'hf87;
      20'h038b7: out <= 12'hb27;
      20'h038b8: out <= 12'hee9;
      20'h038b9: out <= 12'hf87;
      20'h038ba: out <= 12'hee9;
      20'h038bb: out <= 12'hf87;
      20'h038bc: out <= 12'hf87;
      20'h038bd: out <= 12'hb27;
      20'h038be: out <= 12'hf87;
      20'h038bf: out <= 12'hb27;
      20'h038c0: out <= 12'hee9;
      20'h038c1: out <= 12'hf87;
      20'h038c2: out <= 12'hee9;
      20'h038c3: out <= 12'hf87;
      20'h038c4: out <= 12'hf87;
      20'h038c5: out <= 12'hb27;
      20'h038c6: out <= 12'hf87;
      20'h038c7: out <= 12'hb27;
      20'h038c8: out <= 12'hee9;
      20'h038c9: out <= 12'hf87;
      20'h038ca: out <= 12'hee9;
      20'h038cb: out <= 12'hf87;
      20'h038cc: out <= 12'hf87;
      20'h038cd: out <= 12'hb27;
      20'h038ce: out <= 12'hf87;
      20'h038cf: out <= 12'hb27;
      20'h038d0: out <= 12'hee9;
      20'h038d1: out <= 12'hf87;
      20'h038d2: out <= 12'hee9;
      20'h038d3: out <= 12'hf87;
      20'h038d4: out <= 12'hf87;
      20'h038d5: out <= 12'hb27;
      20'h038d6: out <= 12'hf87;
      20'h038d7: out <= 12'hb27;
      20'h038d8: out <= 12'hee9;
      20'h038d9: out <= 12'hf87;
      20'h038da: out <= 12'hee9;
      20'h038db: out <= 12'hf87;
      20'h038dc: out <= 12'hf87;
      20'h038dd: out <= 12'hb27;
      20'h038de: out <= 12'hf87;
      20'h038df: out <= 12'hb27;
      20'h038e0: out <= 12'h000;
      20'h038e1: out <= 12'hfff;
      20'h038e2: out <= 12'hc7f;
      20'h038e3: out <= 12'h72f;
      20'h038e4: out <= 12'hc7f;
      20'h038e5: out <= 12'h72f;
      20'h038e6: out <= 12'h72f;
      20'h038e7: out <= 12'h72f;
      20'h038e8: out <= 12'h72f;
      20'h038e9: out <= 12'h72f;
      20'h038ea: out <= 12'hc7f;
      20'h038eb: out <= 12'hfff;
      20'h038ec: out <= 12'h000;
      20'h038ed: out <= 12'h000;
      20'h038ee: out <= 12'h000;
      20'h038ef: out <= 12'h000;
      20'h038f0: out <= 12'h222;
      20'h038f1: out <= 12'h72f;
      20'h038f2: out <= 12'hc7f;
      20'h038f3: out <= 12'hfff;
      20'h038f4: out <= 12'hc7f;
      20'h038f5: out <= 12'h72f;
      20'h038f6: out <= 12'h72f;
      20'h038f7: out <= 12'h72f;
      20'h038f8: out <= 12'h72f;
      20'h038f9: out <= 12'hfff;
      20'h038fa: out <= 12'hc7f;
      20'h038fb: out <= 12'h72f;
      20'h038fc: out <= 12'h222;
      20'h038fd: out <= 12'h222;
      20'h038fe: out <= 12'h222;
      20'h038ff: out <= 12'h222;
      20'h03900: out <= 12'h000;
      20'h03901: out <= 12'hfff;
      20'h03902: out <= 12'hfff;
      20'h03903: out <= 12'hfff;
      20'h03904: out <= 12'hfff;
      20'h03905: out <= 12'hfff;
      20'h03906: out <= 12'hc7f;
      20'h03907: out <= 12'hc7f;
      20'h03908: out <= 12'hc7f;
      20'h03909: out <= 12'hc7f;
      20'h0390a: out <= 12'hc7f;
      20'h0390b: out <= 12'hfff;
      20'h0390c: out <= 12'hfff;
      20'h0390d: out <= 12'hfff;
      20'h0390e: out <= 12'hfff;
      20'h0390f: out <= 12'hfff;
      20'h03910: out <= 12'h222;
      20'h03911: out <= 12'hfff;
      20'h03912: out <= 12'hfff;
      20'h03913: out <= 12'hfff;
      20'h03914: out <= 12'h72f;
      20'h03915: out <= 12'h72f;
      20'h03916: out <= 12'hc7f;
      20'h03917: out <= 12'hc7f;
      20'h03918: out <= 12'hc7f;
      20'h03919: out <= 12'hc7f;
      20'h0391a: out <= 12'hc7f;
      20'h0391b: out <= 12'h72f;
      20'h0391c: out <= 12'h72f;
      20'h0391d: out <= 12'hfff;
      20'h0391e: out <= 12'hfff;
      20'h0391f: out <= 12'hfff;
      20'h03920: out <= 12'h000;
      20'h03921: out <= 12'h000;
      20'h03922: out <= 12'h000;
      20'h03923: out <= 12'h000;
      20'h03924: out <= 12'hfff;
      20'h03925: out <= 12'hc7f;
      20'h03926: out <= 12'h72f;
      20'h03927: out <= 12'h72f;
      20'h03928: out <= 12'h72f;
      20'h03929: out <= 12'h72f;
      20'h0392a: out <= 12'h72f;
      20'h0392b: out <= 12'hc7f;
      20'h0392c: out <= 12'h72f;
      20'h0392d: out <= 12'hc7f;
      20'h0392e: out <= 12'hfff;
      20'h0392f: out <= 12'h000;
      20'h03930: out <= 12'h222;
      20'h03931: out <= 12'h222;
      20'h03932: out <= 12'h222;
      20'h03933: out <= 12'h222;
      20'h03934: out <= 12'h72f;
      20'h03935: out <= 12'hc7f;
      20'h03936: out <= 12'hfff;
      20'h03937: out <= 12'h72f;
      20'h03938: out <= 12'h72f;
      20'h03939: out <= 12'h72f;
      20'h0393a: out <= 12'h72f;
      20'h0393b: out <= 12'hc7f;
      20'h0393c: out <= 12'hfff;
      20'h0393d: out <= 12'hc7f;
      20'h0393e: out <= 12'h72f;
      20'h0393f: out <= 12'h222;
      20'h03940: out <= 12'h000;
      20'h03941: out <= 12'hfff;
      20'h03942: out <= 12'hc7f;
      20'h03943: out <= 12'h72f;
      20'h03944: out <= 12'h72f;
      20'h03945: out <= 12'hc7f;
      20'h03946: out <= 12'h72f;
      20'h03947: out <= 12'h72f;
      20'h03948: out <= 12'h72f;
      20'h03949: out <= 12'h72f;
      20'h0394a: out <= 12'h72f;
      20'h0394b: out <= 12'hc7f;
      20'h0394c: out <= 12'h72f;
      20'h0394d: out <= 12'h72f;
      20'h0394e: out <= 12'hc7f;
      20'h0394f: out <= 12'hfff;
      20'h03950: out <= 12'h222;
      20'h03951: out <= 12'h72f;
      20'h03952: out <= 12'hc7f;
      20'h03953: out <= 12'hfff;
      20'h03954: out <= 12'h72f;
      20'h03955: out <= 12'hc7f;
      20'h03956: out <= 12'h72f;
      20'h03957: out <= 12'h72f;
      20'h03958: out <= 12'h72f;
      20'h03959: out <= 12'h72f;
      20'h0395a: out <= 12'h72f;
      20'h0395b: out <= 12'hc7f;
      20'h0395c: out <= 12'h72f;
      20'h0395d: out <= 12'hfff;
      20'h0395e: out <= 12'hc7f;
      20'h0395f: out <= 12'h72f;
      20'h03960: out <= 12'h603;
      20'h03961: out <= 12'h603;
      20'h03962: out <= 12'h603;
      20'h03963: out <= 12'h603;
      20'h03964: out <= 12'h000;
      20'h03965: out <= 12'h000;
      20'h03966: out <= 12'hb27;
      20'h03967: out <= 12'hf87;
      20'h03968: out <= 12'hee9;
      20'h03969: out <= 12'hee9;
      20'h0396a: out <= 12'hee9;
      20'h0396b: out <= 12'hee9;
      20'h0396c: out <= 12'hee9;
      20'h0396d: out <= 12'hee9;
      20'h0396e: out <= 12'hee9;
      20'h0396f: out <= 12'hee9;
      20'h03970: out <= 12'hee9;
      20'h03971: out <= 12'hf87;
      20'h03972: out <= 12'hb27;
      20'h03973: out <= 12'h000;
      20'h03974: out <= 12'h000;
      20'h03975: out <= 12'hf87;
      20'h03976: out <= 12'hb27;
      20'h03977: out <= 12'hb27;
      20'h03978: out <= 12'hf87;
      20'h03979: out <= 12'hf87;
      20'h0397a: out <= 12'hf87;
      20'h0397b: out <= 12'hee9;
      20'h0397c: out <= 12'hf87;
      20'h0397d: out <= 12'hee9;
      20'h0397e: out <= 12'hf87;
      20'h0397f: out <= 12'hf87;
      20'h03980: out <= 12'hf87;
      20'h03981: out <= 12'hb27;
      20'h03982: out <= 12'hee9;
      20'h03983: out <= 12'hf87;
      20'h03984: out <= 12'h000;
      20'h03985: out <= 12'h000;
      20'h03986: out <= 12'h000;
      20'h03987: out <= 12'hb27;
      20'h03988: out <= 12'hf87;
      20'h03989: out <= 12'hf87;
      20'h0398a: out <= 12'hf87;
      20'h0398b: out <= 12'hee9;
      20'h0398c: out <= 12'h000;
      20'h0398d: out <= 12'hee9;
      20'h0398e: out <= 12'hf87;
      20'h0398f: out <= 12'h000;
      20'h03990: out <= 12'h000;
      20'h03991: out <= 12'hb27;
      20'h03992: out <= 12'h000;
      20'h03993: out <= 12'hb27;
      20'h03994: out <= 12'h603;
      20'h03995: out <= 12'h603;
      20'h03996: out <= 12'h603;
      20'h03997: out <= 12'h603;
      20'h03998: out <= 12'h603;
      20'h03999: out <= 12'h603;
      20'h0399a: out <= 12'h603;
      20'h0399b: out <= 12'h603;
      20'h0399c: out <= 12'h603;
      20'h0399d: out <= 12'h603;
      20'h0399e: out <= 12'h603;
      20'h0399f: out <= 12'h603;
      20'h039a0: out <= 12'h603;
      20'h039a1: out <= 12'h603;
      20'h039a2: out <= 12'h603;
      20'h039a3: out <= 12'h603;
      20'h039a4: out <= 12'h603;
      20'h039a5: out <= 12'h603;
      20'h039a6: out <= 12'h603;
      20'h039a7: out <= 12'h603;
      20'h039a8: out <= 12'h603;
      20'h039a9: out <= 12'h603;
      20'h039aa: out <= 12'h603;
      20'h039ab: out <= 12'h603;
      20'h039ac: out <= 12'h603;
      20'h039ad: out <= 12'h603;
      20'h039ae: out <= 12'h603;
      20'h039af: out <= 12'h603;
      20'h039b0: out <= 12'h603;
      20'h039b1: out <= 12'h603;
      20'h039b2: out <= 12'h603;
      20'h039b3: out <= 12'h603;
      20'h039b4: out <= 12'h603;
      20'h039b5: out <= 12'h603;
      20'h039b6: out <= 12'h603;
      20'h039b7: out <= 12'h603;
      20'h039b8: out <= 12'hee9;
      20'h039b9: out <= 12'hf87;
      20'h039ba: out <= 12'hee9;
      20'h039bb: out <= 12'hf87;
      20'h039bc: out <= 12'hf87;
      20'h039bd: out <= 12'hb27;
      20'h039be: out <= 12'hf87;
      20'h039bf: out <= 12'hb27;
      20'h039c0: out <= 12'hee9;
      20'h039c1: out <= 12'hf87;
      20'h039c2: out <= 12'hee9;
      20'h039c3: out <= 12'hf87;
      20'h039c4: out <= 12'hf87;
      20'h039c5: out <= 12'hb27;
      20'h039c6: out <= 12'hf87;
      20'h039c7: out <= 12'hb27;
      20'h039c8: out <= 12'hee9;
      20'h039c9: out <= 12'hf87;
      20'h039ca: out <= 12'hee9;
      20'h039cb: out <= 12'hf87;
      20'h039cc: out <= 12'hf87;
      20'h039cd: out <= 12'hb27;
      20'h039ce: out <= 12'hf87;
      20'h039cf: out <= 12'hb27;
      20'h039d0: out <= 12'hee9;
      20'h039d1: out <= 12'hf87;
      20'h039d2: out <= 12'hee9;
      20'h039d3: out <= 12'hf87;
      20'h039d4: out <= 12'hf87;
      20'h039d5: out <= 12'hb27;
      20'h039d6: out <= 12'hf87;
      20'h039d7: out <= 12'hb27;
      20'h039d8: out <= 12'hee9;
      20'h039d9: out <= 12'hf87;
      20'h039da: out <= 12'hee9;
      20'h039db: out <= 12'hf87;
      20'h039dc: out <= 12'hf87;
      20'h039dd: out <= 12'hb27;
      20'h039de: out <= 12'hf87;
      20'h039df: out <= 12'hb27;
      20'h039e0: out <= 12'hee9;
      20'h039e1: out <= 12'hf87;
      20'h039e2: out <= 12'hee9;
      20'h039e3: out <= 12'hf87;
      20'h039e4: out <= 12'hf87;
      20'h039e5: out <= 12'hb27;
      20'h039e6: out <= 12'hf87;
      20'h039e7: out <= 12'hb27;
      20'h039e8: out <= 12'hee9;
      20'h039e9: out <= 12'hf87;
      20'h039ea: out <= 12'hee9;
      20'h039eb: out <= 12'hf87;
      20'h039ec: out <= 12'hf87;
      20'h039ed: out <= 12'hb27;
      20'h039ee: out <= 12'hf87;
      20'h039ef: out <= 12'hb27;
      20'h039f0: out <= 12'hee9;
      20'h039f1: out <= 12'hf87;
      20'h039f2: out <= 12'hee9;
      20'h039f3: out <= 12'hf87;
      20'h039f4: out <= 12'hf87;
      20'h039f5: out <= 12'hb27;
      20'h039f6: out <= 12'hf87;
      20'h039f7: out <= 12'hb27;
      20'h039f8: out <= 12'hfff;
      20'h039f9: out <= 12'hc7f;
      20'h039fa: out <= 12'h72f;
      20'h039fb: out <= 12'hc7f;
      20'h039fc: out <= 12'h72f;
      20'h039fd: out <= 12'h72f;
      20'h039fe: out <= 12'hc7f;
      20'h039ff: out <= 12'hc7f;
      20'h03a00: out <= 12'h72f;
      20'h03a01: out <= 12'h72f;
      20'h03a02: out <= 12'h72f;
      20'h03a03: out <= 12'hc7f;
      20'h03a04: out <= 12'hfff;
      20'h03a05: out <= 12'h000;
      20'h03a06: out <= 12'h000;
      20'h03a07: out <= 12'h000;
      20'h03a08: out <= 12'h72f;
      20'h03a09: out <= 12'hc7f;
      20'h03a0a: out <= 12'hfff;
      20'h03a0b: out <= 12'hc7f;
      20'h03a0c: out <= 12'h72f;
      20'h03a0d: out <= 12'h72f;
      20'h03a0e: out <= 12'hc7f;
      20'h03a0f: out <= 12'hc7f;
      20'h03a10: out <= 12'h72f;
      20'h03a11: out <= 12'h72f;
      20'h03a12: out <= 12'hfff;
      20'h03a13: out <= 12'hc7f;
      20'h03a14: out <= 12'h72f;
      20'h03a15: out <= 12'h222;
      20'h03a16: out <= 12'h222;
      20'h03a17: out <= 12'h222;
      20'h03a18: out <= 12'h000;
      20'h03a19: out <= 12'hc7f;
      20'h03a1a: out <= 12'h72f;
      20'h03a1b: out <= 12'hfff;
      20'h03a1c: out <= 12'hc7f;
      20'h03a1d: out <= 12'hc7f;
      20'h03a1e: out <= 12'h72f;
      20'h03a1f: out <= 12'h72f;
      20'h03a20: out <= 12'h72f;
      20'h03a21: out <= 12'h72f;
      20'h03a22: out <= 12'h72f;
      20'h03a23: out <= 12'hc7f;
      20'h03a24: out <= 12'hc7f;
      20'h03a25: out <= 12'hfff;
      20'h03a26: out <= 12'h72f;
      20'h03a27: out <= 12'hc7f;
      20'h03a28: out <= 12'h222;
      20'h03a29: out <= 12'hc7f;
      20'h03a2a: out <= 12'h72f;
      20'h03a2b: out <= 12'h72f;
      20'h03a2c: out <= 12'hc7f;
      20'h03a2d: out <= 12'hc7f;
      20'h03a2e: out <= 12'hfff;
      20'h03a2f: out <= 12'hfff;
      20'h03a30: out <= 12'hfff;
      20'h03a31: out <= 12'hfff;
      20'h03a32: out <= 12'hfff;
      20'h03a33: out <= 12'hc7f;
      20'h03a34: out <= 12'hc7f;
      20'h03a35: out <= 12'h72f;
      20'h03a36: out <= 12'h72f;
      20'h03a37: out <= 12'hc7f;
      20'h03a38: out <= 12'h000;
      20'h03a39: out <= 12'h000;
      20'h03a3a: out <= 12'h000;
      20'h03a3b: out <= 12'hfff;
      20'h03a3c: out <= 12'hc7f;
      20'h03a3d: out <= 12'h72f;
      20'h03a3e: out <= 12'h72f;
      20'h03a3f: out <= 12'h72f;
      20'h03a40: out <= 12'hc7f;
      20'h03a41: out <= 12'hc7f;
      20'h03a42: out <= 12'h72f;
      20'h03a43: out <= 12'h72f;
      20'h03a44: out <= 12'hc7f;
      20'h03a45: out <= 12'h72f;
      20'h03a46: out <= 12'hc7f;
      20'h03a47: out <= 12'hfff;
      20'h03a48: out <= 12'h222;
      20'h03a49: out <= 12'h222;
      20'h03a4a: out <= 12'h222;
      20'h03a4b: out <= 12'h72f;
      20'h03a4c: out <= 12'hc7f;
      20'h03a4d: out <= 12'hfff;
      20'h03a4e: out <= 12'h72f;
      20'h03a4f: out <= 12'h72f;
      20'h03a50: out <= 12'hc7f;
      20'h03a51: out <= 12'hc7f;
      20'h03a52: out <= 12'h72f;
      20'h03a53: out <= 12'h72f;
      20'h03a54: out <= 12'hc7f;
      20'h03a55: out <= 12'hfff;
      20'h03a56: out <= 12'hc7f;
      20'h03a57: out <= 12'h72f;
      20'h03a58: out <= 12'h000;
      20'h03a59: out <= 12'hfff;
      20'h03a5a: out <= 12'hc7f;
      20'h03a5b: out <= 12'h72f;
      20'h03a5c: out <= 12'h72f;
      20'h03a5d: out <= 12'h72f;
      20'h03a5e: out <= 12'h72f;
      20'h03a5f: out <= 12'hc7f;
      20'h03a60: out <= 12'hfff;
      20'h03a61: out <= 12'hc7f;
      20'h03a62: out <= 12'h72f;
      20'h03a63: out <= 12'h72f;
      20'h03a64: out <= 12'h72f;
      20'h03a65: out <= 12'h72f;
      20'h03a66: out <= 12'hc7f;
      20'h03a67: out <= 12'hfff;
      20'h03a68: out <= 12'h222;
      20'h03a69: out <= 12'h72f;
      20'h03a6a: out <= 12'hc7f;
      20'h03a6b: out <= 12'hfff;
      20'h03a6c: out <= 12'h72f;
      20'h03a6d: out <= 12'h72f;
      20'h03a6e: out <= 12'h72f;
      20'h03a6f: out <= 12'hc7f;
      20'h03a70: out <= 12'hfff;
      20'h03a71: out <= 12'hc7f;
      20'h03a72: out <= 12'h72f;
      20'h03a73: out <= 12'h72f;
      20'h03a74: out <= 12'h72f;
      20'h03a75: out <= 12'hfff;
      20'h03a76: out <= 12'hc7f;
      20'h03a77: out <= 12'h72f;
      20'h03a78: out <= 12'h603;
      20'h03a79: out <= 12'h603;
      20'h03a7a: out <= 12'h603;
      20'h03a7b: out <= 12'h603;
      20'h03a7c: out <= 12'h000;
      20'h03a7d: out <= 12'h000;
      20'h03a7e: out <= 12'hb27;
      20'h03a7f: out <= 12'hf87;
      20'h03a80: out <= 12'hee9;
      20'h03a81: out <= 12'hee9;
      20'h03a82: out <= 12'hee9;
      20'h03a83: out <= 12'hee9;
      20'h03a84: out <= 12'hee9;
      20'h03a85: out <= 12'hee9;
      20'h03a86: out <= 12'hee9;
      20'h03a87: out <= 12'hee9;
      20'h03a88: out <= 12'hee9;
      20'h03a89: out <= 12'hf87;
      20'h03a8a: out <= 12'hb27;
      20'h03a8b: out <= 12'h000;
      20'h03a8c: out <= 12'h000;
      20'h03a8d: out <= 12'hf87;
      20'h03a8e: out <= 12'hb27;
      20'h03a8f: out <= 12'hf87;
      20'h03a90: out <= 12'hb27;
      20'h03a91: out <= 12'hf87;
      20'h03a92: out <= 12'hf87;
      20'h03a93: out <= 12'hf87;
      20'h03a94: out <= 12'hee9;
      20'h03a95: out <= 12'hf87;
      20'h03a96: out <= 12'hf87;
      20'h03a97: out <= 12'hf87;
      20'h03a98: out <= 12'hb27;
      20'h03a99: out <= 12'hf87;
      20'h03a9a: out <= 12'hee9;
      20'h03a9b: out <= 12'hf87;
      20'h03a9c: out <= 12'h000;
      20'h03a9d: out <= 12'h000;
      20'h03a9e: out <= 12'h000;
      20'h03a9f: out <= 12'h000;
      20'h03aa0: out <= 12'hb27;
      20'h03aa1: out <= 12'hf87;
      20'h03aa2: out <= 12'hf87;
      20'h03aa3: out <= 12'hf87;
      20'h03aa4: out <= 12'hee9;
      20'h03aa5: out <= 12'hf87;
      20'h03aa6: out <= 12'hf87;
      20'h03aa7: out <= 12'hf87;
      20'h03aa8: out <= 12'hb27;
      20'h03aa9: out <= 12'h000;
      20'h03aaa: out <= 12'hb27;
      20'h03aab: out <= 12'hb27;
      20'h03aac: out <= 12'h603;
      20'h03aad: out <= 12'h603;
      20'h03aae: out <= 12'h603;
      20'h03aaf: out <= 12'h603;
      20'h03ab0: out <= 12'h603;
      20'h03ab1: out <= 12'h603;
      20'h03ab2: out <= 12'h603;
      20'h03ab3: out <= 12'h603;
      20'h03ab4: out <= 12'h603;
      20'h03ab5: out <= 12'h603;
      20'h03ab6: out <= 12'h603;
      20'h03ab7: out <= 12'h603;
      20'h03ab8: out <= 12'h603;
      20'h03ab9: out <= 12'h603;
      20'h03aba: out <= 12'h603;
      20'h03abb: out <= 12'h603;
      20'h03abc: out <= 12'h603;
      20'h03abd: out <= 12'h603;
      20'h03abe: out <= 12'h603;
      20'h03abf: out <= 12'h603;
      20'h03ac0: out <= 12'h603;
      20'h03ac1: out <= 12'h603;
      20'h03ac2: out <= 12'h603;
      20'h03ac3: out <= 12'h603;
      20'h03ac4: out <= 12'h603;
      20'h03ac5: out <= 12'h603;
      20'h03ac6: out <= 12'h603;
      20'h03ac7: out <= 12'h603;
      20'h03ac8: out <= 12'h603;
      20'h03ac9: out <= 12'h603;
      20'h03aca: out <= 12'h603;
      20'h03acb: out <= 12'h603;
      20'h03acc: out <= 12'h603;
      20'h03acd: out <= 12'h603;
      20'h03ace: out <= 12'h603;
      20'h03acf: out <= 12'h603;
      20'h03ad0: out <= 12'hee9;
      20'h03ad1: out <= 12'hf87;
      20'h03ad2: out <= 12'hee9;
      20'h03ad3: out <= 12'hb27;
      20'h03ad4: out <= 12'hb27;
      20'h03ad5: out <= 12'hb27;
      20'h03ad6: out <= 12'hf87;
      20'h03ad7: out <= 12'hb27;
      20'h03ad8: out <= 12'hee9;
      20'h03ad9: out <= 12'hf87;
      20'h03ada: out <= 12'hee9;
      20'h03adb: out <= 12'hb27;
      20'h03adc: out <= 12'hb27;
      20'h03add: out <= 12'hb27;
      20'h03ade: out <= 12'hf87;
      20'h03adf: out <= 12'hb27;
      20'h03ae0: out <= 12'hee9;
      20'h03ae1: out <= 12'hf87;
      20'h03ae2: out <= 12'hee9;
      20'h03ae3: out <= 12'hb27;
      20'h03ae4: out <= 12'hb27;
      20'h03ae5: out <= 12'hb27;
      20'h03ae6: out <= 12'hf87;
      20'h03ae7: out <= 12'hb27;
      20'h03ae8: out <= 12'hee9;
      20'h03ae9: out <= 12'hf87;
      20'h03aea: out <= 12'hee9;
      20'h03aeb: out <= 12'hb27;
      20'h03aec: out <= 12'hb27;
      20'h03aed: out <= 12'hb27;
      20'h03aee: out <= 12'hf87;
      20'h03aef: out <= 12'hb27;
      20'h03af0: out <= 12'hee9;
      20'h03af1: out <= 12'hf87;
      20'h03af2: out <= 12'hee9;
      20'h03af3: out <= 12'hb27;
      20'h03af4: out <= 12'hb27;
      20'h03af5: out <= 12'hb27;
      20'h03af6: out <= 12'hf87;
      20'h03af7: out <= 12'hb27;
      20'h03af8: out <= 12'hee9;
      20'h03af9: out <= 12'hf87;
      20'h03afa: out <= 12'hee9;
      20'h03afb: out <= 12'hb27;
      20'h03afc: out <= 12'hb27;
      20'h03afd: out <= 12'hb27;
      20'h03afe: out <= 12'hf87;
      20'h03aff: out <= 12'hb27;
      20'h03b00: out <= 12'hee9;
      20'h03b01: out <= 12'hf87;
      20'h03b02: out <= 12'hee9;
      20'h03b03: out <= 12'hb27;
      20'h03b04: out <= 12'hb27;
      20'h03b05: out <= 12'hb27;
      20'h03b06: out <= 12'hf87;
      20'h03b07: out <= 12'hb27;
      20'h03b08: out <= 12'hee9;
      20'h03b09: out <= 12'hf87;
      20'h03b0a: out <= 12'hee9;
      20'h03b0b: out <= 12'hb27;
      20'h03b0c: out <= 12'hb27;
      20'h03b0d: out <= 12'hb27;
      20'h03b0e: out <= 12'hf87;
      20'h03b0f: out <= 12'hb27;
      20'h03b10: out <= 12'hfff;
      20'h03b11: out <= 12'hc7f;
      20'h03b12: out <= 12'h72f;
      20'h03b13: out <= 12'hfff;
      20'h03b14: out <= 12'h72f;
      20'h03b15: out <= 12'hc7f;
      20'h03b16: out <= 12'hfff;
      20'h03b17: out <= 12'hfff;
      20'h03b18: out <= 12'hc7f;
      20'h03b19: out <= 12'h72f;
      20'h03b1a: out <= 12'h72f;
      20'h03b1b: out <= 12'hc7f;
      20'h03b1c: out <= 12'hfff;
      20'h03b1d: out <= 12'h72f;
      20'h03b1e: out <= 12'h72f;
      20'h03b1f: out <= 12'hc7f;
      20'h03b20: out <= 12'h72f;
      20'h03b21: out <= 12'hc7f;
      20'h03b22: out <= 12'hfff;
      20'h03b23: out <= 12'hfff;
      20'h03b24: out <= 12'h72f;
      20'h03b25: out <= 12'hc7f;
      20'h03b26: out <= 12'hfff;
      20'h03b27: out <= 12'hfff;
      20'h03b28: out <= 12'hc7f;
      20'h03b29: out <= 12'h72f;
      20'h03b2a: out <= 12'hfff;
      20'h03b2b: out <= 12'hc7f;
      20'h03b2c: out <= 12'h72f;
      20'h03b2d: out <= 12'h72f;
      20'h03b2e: out <= 12'h72f;
      20'h03b2f: out <= 12'hc7f;
      20'h03b30: out <= 12'h000;
      20'h03b31: out <= 12'hc7f;
      20'h03b32: out <= 12'hfff;
      20'h03b33: out <= 12'hc7f;
      20'h03b34: out <= 12'h72f;
      20'h03b35: out <= 12'h72f;
      20'h03b36: out <= 12'h72f;
      20'h03b37: out <= 12'h72f;
      20'h03b38: out <= 12'h72f;
      20'h03b39: out <= 12'h72f;
      20'h03b3a: out <= 12'h72f;
      20'h03b3b: out <= 12'h72f;
      20'h03b3c: out <= 12'h72f;
      20'h03b3d: out <= 12'hc7f;
      20'h03b3e: out <= 12'hfff;
      20'h03b3f: out <= 12'hc7f;
      20'h03b40: out <= 12'h222;
      20'h03b41: out <= 12'hc7f;
      20'h03b42: out <= 12'h72f;
      20'h03b43: out <= 12'hc7f;
      20'h03b44: out <= 12'hfff;
      20'h03b45: out <= 12'hfff;
      20'h03b46: out <= 12'h72f;
      20'h03b47: out <= 12'h72f;
      20'h03b48: out <= 12'h72f;
      20'h03b49: out <= 12'h72f;
      20'h03b4a: out <= 12'h72f;
      20'h03b4b: out <= 12'hfff;
      20'h03b4c: out <= 12'hfff;
      20'h03b4d: out <= 12'hc7f;
      20'h03b4e: out <= 12'h72f;
      20'h03b4f: out <= 12'hc7f;
      20'h03b50: out <= 12'hc7f;
      20'h03b51: out <= 12'h72f;
      20'h03b52: out <= 12'h72f;
      20'h03b53: out <= 12'hfff;
      20'h03b54: out <= 12'hc7f;
      20'h03b55: out <= 12'h72f;
      20'h03b56: out <= 12'h72f;
      20'h03b57: out <= 12'hc7f;
      20'h03b58: out <= 12'hfff;
      20'h03b59: out <= 12'hfff;
      20'h03b5a: out <= 12'hc7f;
      20'h03b5b: out <= 12'h72f;
      20'h03b5c: out <= 12'hfff;
      20'h03b5d: out <= 12'h72f;
      20'h03b5e: out <= 12'hc7f;
      20'h03b5f: out <= 12'hfff;
      20'h03b60: out <= 12'hc7f;
      20'h03b61: out <= 12'h72f;
      20'h03b62: out <= 12'h72f;
      20'h03b63: out <= 12'h72f;
      20'h03b64: out <= 12'hc7f;
      20'h03b65: out <= 12'hfff;
      20'h03b66: out <= 12'h72f;
      20'h03b67: out <= 12'hc7f;
      20'h03b68: out <= 12'hfff;
      20'h03b69: out <= 12'hfff;
      20'h03b6a: out <= 12'hc7f;
      20'h03b6b: out <= 12'h72f;
      20'h03b6c: out <= 12'hfff;
      20'h03b6d: out <= 12'hfff;
      20'h03b6e: out <= 12'hc7f;
      20'h03b6f: out <= 12'h72f;
      20'h03b70: out <= 12'h000;
      20'h03b71: out <= 12'hfff;
      20'h03b72: out <= 12'hc7f;
      20'h03b73: out <= 12'h72f;
      20'h03b74: out <= 12'h72f;
      20'h03b75: out <= 12'h72f;
      20'h03b76: out <= 12'hc7f;
      20'h03b77: out <= 12'hfff;
      20'h03b78: out <= 12'hfff;
      20'h03b79: out <= 12'hfff;
      20'h03b7a: out <= 12'hc7f;
      20'h03b7b: out <= 12'h72f;
      20'h03b7c: out <= 12'h72f;
      20'h03b7d: out <= 12'h72f;
      20'h03b7e: out <= 12'hc7f;
      20'h03b7f: out <= 12'hfff;
      20'h03b80: out <= 12'h222;
      20'h03b81: out <= 12'h72f;
      20'h03b82: out <= 12'hc7f;
      20'h03b83: out <= 12'hfff;
      20'h03b84: out <= 12'h72f;
      20'h03b85: out <= 12'h72f;
      20'h03b86: out <= 12'hc7f;
      20'h03b87: out <= 12'hfff;
      20'h03b88: out <= 12'hfff;
      20'h03b89: out <= 12'hfff;
      20'h03b8a: out <= 12'hc7f;
      20'h03b8b: out <= 12'h72f;
      20'h03b8c: out <= 12'h72f;
      20'h03b8d: out <= 12'hfff;
      20'h03b8e: out <= 12'hc7f;
      20'h03b8f: out <= 12'h72f;
      20'h03b90: out <= 12'h603;
      20'h03b91: out <= 12'h603;
      20'h03b92: out <= 12'h603;
      20'h03b93: out <= 12'h603;
      20'h03b94: out <= 12'h000;
      20'h03b95: out <= 12'h000;
      20'h03b96: out <= 12'hb27;
      20'h03b97: out <= 12'hf87;
      20'h03b98: out <= 12'hee9;
      20'h03b99: out <= 12'hee9;
      20'h03b9a: out <= 12'hee9;
      20'h03b9b: out <= 12'hee9;
      20'h03b9c: out <= 12'hee9;
      20'h03b9d: out <= 12'hee9;
      20'h03b9e: out <= 12'hee9;
      20'h03b9f: out <= 12'hee9;
      20'h03ba0: out <= 12'hf87;
      20'h03ba1: out <= 12'hf87;
      20'h03ba2: out <= 12'hb27;
      20'h03ba3: out <= 12'h000;
      20'h03ba4: out <= 12'h000;
      20'h03ba5: out <= 12'hf87;
      20'h03ba6: out <= 12'hb27;
      20'h03ba7: out <= 12'hf87;
      20'h03ba8: out <= 12'hf87;
      20'h03ba9: out <= 12'hb27;
      20'h03baa: out <= 12'hf87;
      20'h03bab: out <= 12'hee9;
      20'h03bac: out <= 12'hf87;
      20'h03bad: out <= 12'hf87;
      20'h03bae: out <= 12'hf87;
      20'h03baf: out <= 12'hb27;
      20'h03bb0: out <= 12'hf87;
      20'h03bb1: out <= 12'hf87;
      20'h03bb2: out <= 12'hee9;
      20'h03bb3: out <= 12'hf87;
      20'h03bb4: out <= 12'h000;
      20'h03bb5: out <= 12'h000;
      20'h03bb6: out <= 12'h000;
      20'h03bb7: out <= 12'h000;
      20'h03bb8: out <= 12'h000;
      20'h03bb9: out <= 12'hb27;
      20'h03bba: out <= 12'hf87;
      20'h03bbb: out <= 12'hee9;
      20'h03bbc: out <= 12'hf87;
      20'h03bbd: out <= 12'hf87;
      20'h03bbe: out <= 12'hf87;
      20'h03bbf: out <= 12'hb27;
      20'h03bc0: out <= 12'hb27;
      20'h03bc1: out <= 12'hb27;
      20'h03bc2: out <= 12'hb27;
      20'h03bc3: out <= 12'hb27;
      20'h03bc4: out <= 12'h603;
      20'h03bc5: out <= 12'h603;
      20'h03bc6: out <= 12'h603;
      20'h03bc7: out <= 12'h603;
      20'h03bc8: out <= 12'h603;
      20'h03bc9: out <= 12'h603;
      20'h03bca: out <= 12'h603;
      20'h03bcb: out <= 12'h603;
      20'h03bcc: out <= 12'h603;
      20'h03bcd: out <= 12'h603;
      20'h03bce: out <= 12'h603;
      20'h03bcf: out <= 12'h603;
      20'h03bd0: out <= 12'h603;
      20'h03bd1: out <= 12'h603;
      20'h03bd2: out <= 12'h603;
      20'h03bd3: out <= 12'h603;
      20'h03bd4: out <= 12'h603;
      20'h03bd5: out <= 12'h603;
      20'h03bd6: out <= 12'h603;
      20'h03bd7: out <= 12'h603;
      20'h03bd8: out <= 12'h603;
      20'h03bd9: out <= 12'h603;
      20'h03bda: out <= 12'h603;
      20'h03bdb: out <= 12'h603;
      20'h03bdc: out <= 12'h603;
      20'h03bdd: out <= 12'h603;
      20'h03bde: out <= 12'h603;
      20'h03bdf: out <= 12'h603;
      20'h03be0: out <= 12'h603;
      20'h03be1: out <= 12'h603;
      20'h03be2: out <= 12'h603;
      20'h03be3: out <= 12'h603;
      20'h03be4: out <= 12'h603;
      20'h03be5: out <= 12'h603;
      20'h03be6: out <= 12'h603;
      20'h03be7: out <= 12'h603;
      20'h03be8: out <= 12'hee9;
      20'h03be9: out <= 12'hf87;
      20'h03bea: out <= 12'hf87;
      20'h03beb: out <= 12'hf87;
      20'h03bec: out <= 12'hf87;
      20'h03bed: out <= 12'hf87;
      20'h03bee: out <= 12'hf87;
      20'h03bef: out <= 12'hb27;
      20'h03bf0: out <= 12'hee9;
      20'h03bf1: out <= 12'hf87;
      20'h03bf2: out <= 12'hf87;
      20'h03bf3: out <= 12'hf87;
      20'h03bf4: out <= 12'hf87;
      20'h03bf5: out <= 12'hf87;
      20'h03bf6: out <= 12'hf87;
      20'h03bf7: out <= 12'hb27;
      20'h03bf8: out <= 12'hee9;
      20'h03bf9: out <= 12'hf87;
      20'h03bfa: out <= 12'hf87;
      20'h03bfb: out <= 12'hf87;
      20'h03bfc: out <= 12'hf87;
      20'h03bfd: out <= 12'hf87;
      20'h03bfe: out <= 12'hf87;
      20'h03bff: out <= 12'hb27;
      20'h03c00: out <= 12'hee9;
      20'h03c01: out <= 12'hf87;
      20'h03c02: out <= 12'hf87;
      20'h03c03: out <= 12'hf87;
      20'h03c04: out <= 12'hf87;
      20'h03c05: out <= 12'hf87;
      20'h03c06: out <= 12'hf87;
      20'h03c07: out <= 12'hb27;
      20'h03c08: out <= 12'hee9;
      20'h03c09: out <= 12'hf87;
      20'h03c0a: out <= 12'hf87;
      20'h03c0b: out <= 12'hf87;
      20'h03c0c: out <= 12'hf87;
      20'h03c0d: out <= 12'hf87;
      20'h03c0e: out <= 12'hf87;
      20'h03c0f: out <= 12'hb27;
      20'h03c10: out <= 12'hee9;
      20'h03c11: out <= 12'hf87;
      20'h03c12: out <= 12'hf87;
      20'h03c13: out <= 12'hf87;
      20'h03c14: out <= 12'hf87;
      20'h03c15: out <= 12'hf87;
      20'h03c16: out <= 12'hf87;
      20'h03c17: out <= 12'hb27;
      20'h03c18: out <= 12'hee9;
      20'h03c19: out <= 12'hf87;
      20'h03c1a: out <= 12'hf87;
      20'h03c1b: out <= 12'hf87;
      20'h03c1c: out <= 12'hf87;
      20'h03c1d: out <= 12'hf87;
      20'h03c1e: out <= 12'hf87;
      20'h03c1f: out <= 12'hb27;
      20'h03c20: out <= 12'hee9;
      20'h03c21: out <= 12'hf87;
      20'h03c22: out <= 12'hf87;
      20'h03c23: out <= 12'hf87;
      20'h03c24: out <= 12'hf87;
      20'h03c25: out <= 12'hf87;
      20'h03c26: out <= 12'hf87;
      20'h03c27: out <= 12'hb27;
      20'h03c28: out <= 12'hfff;
      20'h03c29: out <= 12'hc7f;
      20'h03c2a: out <= 12'h72f;
      20'h03c2b: out <= 12'hfff;
      20'h03c2c: out <= 12'h72f;
      20'h03c2d: out <= 12'hfff;
      20'h03c2e: out <= 12'hfff;
      20'h03c2f: out <= 12'hfff;
      20'h03c30: out <= 12'hfff;
      20'h03c31: out <= 12'h72f;
      20'h03c32: out <= 12'h72f;
      20'h03c33: out <= 12'hc7f;
      20'h03c34: out <= 12'hfff;
      20'h03c35: out <= 12'hfff;
      20'h03c36: out <= 12'hfff;
      20'h03c37: out <= 12'hfff;
      20'h03c38: out <= 12'h72f;
      20'h03c39: out <= 12'hc7f;
      20'h03c3a: out <= 12'hfff;
      20'h03c3b: out <= 12'hfff;
      20'h03c3c: out <= 12'h72f;
      20'h03c3d: out <= 12'hfff;
      20'h03c3e: out <= 12'hfff;
      20'h03c3f: out <= 12'hfff;
      20'h03c40: out <= 12'hfff;
      20'h03c41: out <= 12'h72f;
      20'h03c42: out <= 12'hfff;
      20'h03c43: out <= 12'hc7f;
      20'h03c44: out <= 12'h72f;
      20'h03c45: out <= 12'hfff;
      20'h03c46: out <= 12'hfff;
      20'h03c47: out <= 12'hfff;
      20'h03c48: out <= 12'h000;
      20'h03c49: out <= 12'hfff;
      20'h03c4a: out <= 12'hc7f;
      20'h03c4b: out <= 12'h72f;
      20'h03c4c: out <= 12'h72f;
      20'h03c4d: out <= 12'h72f;
      20'h03c4e: out <= 12'h72f;
      20'h03c4f: out <= 12'hc7f;
      20'h03c50: out <= 12'hfff;
      20'h03c51: out <= 12'hc7f;
      20'h03c52: out <= 12'h72f;
      20'h03c53: out <= 12'h72f;
      20'h03c54: out <= 12'h72f;
      20'h03c55: out <= 12'h72f;
      20'h03c56: out <= 12'hc7f;
      20'h03c57: out <= 12'hfff;
      20'h03c58: out <= 12'h222;
      20'h03c59: out <= 12'h72f;
      20'h03c5a: out <= 12'hc7f;
      20'h03c5b: out <= 12'hfff;
      20'h03c5c: out <= 12'h72f;
      20'h03c5d: out <= 12'h72f;
      20'h03c5e: out <= 12'h72f;
      20'h03c5f: out <= 12'hc7f;
      20'h03c60: out <= 12'hfff;
      20'h03c61: out <= 12'hc7f;
      20'h03c62: out <= 12'h72f;
      20'h03c63: out <= 12'h72f;
      20'h03c64: out <= 12'h72f;
      20'h03c65: out <= 12'hfff;
      20'h03c66: out <= 12'hc7f;
      20'h03c67: out <= 12'h72f;
      20'h03c68: out <= 12'hfff;
      20'h03c69: out <= 12'hfff;
      20'h03c6a: out <= 12'hfff;
      20'h03c6b: out <= 12'hfff;
      20'h03c6c: out <= 12'hc7f;
      20'h03c6d: out <= 12'h72f;
      20'h03c6e: out <= 12'h72f;
      20'h03c6f: out <= 12'hfff;
      20'h03c70: out <= 12'hfff;
      20'h03c71: out <= 12'hfff;
      20'h03c72: out <= 12'hfff;
      20'h03c73: out <= 12'h72f;
      20'h03c74: out <= 12'hfff;
      20'h03c75: out <= 12'h72f;
      20'h03c76: out <= 12'hc7f;
      20'h03c77: out <= 12'hfff;
      20'h03c78: out <= 12'hfff;
      20'h03c79: out <= 12'hfff;
      20'h03c7a: out <= 12'hfff;
      20'h03c7b: out <= 12'h72f;
      20'h03c7c: out <= 12'hc7f;
      20'h03c7d: out <= 12'hfff;
      20'h03c7e: out <= 12'h72f;
      20'h03c7f: out <= 12'hfff;
      20'h03c80: out <= 12'hfff;
      20'h03c81: out <= 12'hfff;
      20'h03c82: out <= 12'hfff;
      20'h03c83: out <= 12'h72f;
      20'h03c84: out <= 12'hfff;
      20'h03c85: out <= 12'hfff;
      20'h03c86: out <= 12'hc7f;
      20'h03c87: out <= 12'h72f;
      20'h03c88: out <= 12'h000;
      20'h03c89: out <= 12'hfff;
      20'h03c8a: out <= 12'hc7f;
      20'h03c8b: out <= 12'h72f;
      20'h03c8c: out <= 12'h72f;
      20'h03c8d: out <= 12'h72f;
      20'h03c8e: out <= 12'hc7f;
      20'h03c8f: out <= 12'hfff;
      20'h03c90: out <= 12'hfff;
      20'h03c91: out <= 12'hfff;
      20'h03c92: out <= 12'hc7f;
      20'h03c93: out <= 12'h72f;
      20'h03c94: out <= 12'h72f;
      20'h03c95: out <= 12'h72f;
      20'h03c96: out <= 12'hc7f;
      20'h03c97: out <= 12'hfff;
      20'h03c98: out <= 12'h222;
      20'h03c99: out <= 12'h72f;
      20'h03c9a: out <= 12'hc7f;
      20'h03c9b: out <= 12'hfff;
      20'h03c9c: out <= 12'h72f;
      20'h03c9d: out <= 12'h72f;
      20'h03c9e: out <= 12'hc7f;
      20'h03c9f: out <= 12'hfff;
      20'h03ca0: out <= 12'hfff;
      20'h03ca1: out <= 12'hfff;
      20'h03ca2: out <= 12'hc7f;
      20'h03ca3: out <= 12'h72f;
      20'h03ca4: out <= 12'h72f;
      20'h03ca5: out <= 12'hfff;
      20'h03ca6: out <= 12'hc7f;
      20'h03ca7: out <= 12'h72f;
      20'h03ca8: out <= 12'h603;
      20'h03ca9: out <= 12'h603;
      20'h03caa: out <= 12'h603;
      20'h03cab: out <= 12'h603;
      20'h03cac: out <= 12'h000;
      20'h03cad: out <= 12'h000;
      20'h03cae: out <= 12'hb27;
      20'h03caf: out <= 12'hf87;
      20'h03cb0: out <= 12'hee9;
      20'h03cb1: out <= 12'hee9;
      20'h03cb2: out <= 12'hee9;
      20'h03cb3: out <= 12'hee9;
      20'h03cb4: out <= 12'hee9;
      20'h03cb5: out <= 12'hee9;
      20'h03cb6: out <= 12'hee9;
      20'h03cb7: out <= 12'hf87;
      20'h03cb8: out <= 12'hee9;
      20'h03cb9: out <= 12'hf87;
      20'h03cba: out <= 12'hb27;
      20'h03cbb: out <= 12'h000;
      20'h03cbc: out <= 12'h000;
      20'h03cbd: out <= 12'hf87;
      20'h03cbe: out <= 12'hb27;
      20'h03cbf: out <= 12'hf87;
      20'h03cc0: out <= 12'hf87;
      20'h03cc1: out <= 12'hf87;
      20'h03cc2: out <= 12'hee9;
      20'h03cc3: out <= 12'hf87;
      20'h03cc4: out <= 12'hf87;
      20'h03cc5: out <= 12'hf87;
      20'h03cc6: out <= 12'hb27;
      20'h03cc7: out <= 12'hf87;
      20'h03cc8: out <= 12'hf87;
      20'h03cc9: out <= 12'hf87;
      20'h03cca: out <= 12'hee9;
      20'h03ccb: out <= 12'hf87;
      20'h03ccc: out <= 12'h000;
      20'h03ccd: out <= 12'h000;
      20'h03cce: out <= 12'h000;
      20'h03ccf: out <= 12'hb27;
      20'h03cd0: out <= 12'h000;
      20'h03cd1: out <= 12'hb27;
      20'h03cd2: out <= 12'hee9;
      20'h03cd3: out <= 12'hf87;
      20'h03cd4: out <= 12'hf87;
      20'h03cd5: out <= 12'hf87;
      20'h03cd6: out <= 12'hb27;
      20'h03cd7: out <= 12'hf87;
      20'h03cd8: out <= 12'hb27;
      20'h03cd9: out <= 12'hb27;
      20'h03cda: out <= 12'hb27;
      20'h03cdb: out <= 12'hf87;
      20'h03cdc: out <= 12'h603;
      20'h03cdd: out <= 12'h603;
      20'h03cde: out <= 12'h603;
      20'h03cdf: out <= 12'h603;
      20'h03ce0: out <= 12'h603;
      20'h03ce1: out <= 12'h603;
      20'h03ce2: out <= 12'h603;
      20'h03ce3: out <= 12'h603;
      20'h03ce4: out <= 12'h603;
      20'h03ce5: out <= 12'h603;
      20'h03ce6: out <= 12'h603;
      20'h03ce7: out <= 12'h603;
      20'h03ce8: out <= 12'h603;
      20'h03ce9: out <= 12'h603;
      20'h03cea: out <= 12'h603;
      20'h03ceb: out <= 12'h603;
      20'h03cec: out <= 12'h603;
      20'h03ced: out <= 12'h603;
      20'h03cee: out <= 12'h603;
      20'h03cef: out <= 12'h603;
      20'h03cf0: out <= 12'h603;
      20'h03cf1: out <= 12'h603;
      20'h03cf2: out <= 12'h603;
      20'h03cf3: out <= 12'h603;
      20'h03cf4: out <= 12'h603;
      20'h03cf5: out <= 12'h603;
      20'h03cf6: out <= 12'h603;
      20'h03cf7: out <= 12'h603;
      20'h03cf8: out <= 12'h603;
      20'h03cf9: out <= 12'h603;
      20'h03cfa: out <= 12'h603;
      20'h03cfb: out <= 12'h603;
      20'h03cfc: out <= 12'h603;
      20'h03cfd: out <= 12'h603;
      20'h03cfe: out <= 12'h603;
      20'h03cff: out <= 12'h603;
      20'h03d00: out <= 12'hb27;
      20'h03d01: out <= 12'hb27;
      20'h03d02: out <= 12'hb27;
      20'h03d03: out <= 12'hb27;
      20'h03d04: out <= 12'hb27;
      20'h03d05: out <= 12'hb27;
      20'h03d06: out <= 12'hb27;
      20'h03d07: out <= 12'hb27;
      20'h03d08: out <= 12'hb27;
      20'h03d09: out <= 12'hb27;
      20'h03d0a: out <= 12'hb27;
      20'h03d0b: out <= 12'hb27;
      20'h03d0c: out <= 12'hb27;
      20'h03d0d: out <= 12'hb27;
      20'h03d0e: out <= 12'hb27;
      20'h03d0f: out <= 12'hb27;
      20'h03d10: out <= 12'hb27;
      20'h03d11: out <= 12'hb27;
      20'h03d12: out <= 12'hb27;
      20'h03d13: out <= 12'hb27;
      20'h03d14: out <= 12'hb27;
      20'h03d15: out <= 12'hb27;
      20'h03d16: out <= 12'hb27;
      20'h03d17: out <= 12'hb27;
      20'h03d18: out <= 12'hb27;
      20'h03d19: out <= 12'hb27;
      20'h03d1a: out <= 12'hb27;
      20'h03d1b: out <= 12'hb27;
      20'h03d1c: out <= 12'hb27;
      20'h03d1d: out <= 12'hb27;
      20'h03d1e: out <= 12'hb27;
      20'h03d1f: out <= 12'hb27;
      20'h03d20: out <= 12'hb27;
      20'h03d21: out <= 12'hb27;
      20'h03d22: out <= 12'hb27;
      20'h03d23: out <= 12'hb27;
      20'h03d24: out <= 12'hb27;
      20'h03d25: out <= 12'hb27;
      20'h03d26: out <= 12'hb27;
      20'h03d27: out <= 12'hb27;
      20'h03d28: out <= 12'hb27;
      20'h03d29: out <= 12'hb27;
      20'h03d2a: out <= 12'hb27;
      20'h03d2b: out <= 12'hb27;
      20'h03d2c: out <= 12'hb27;
      20'h03d2d: out <= 12'hb27;
      20'h03d2e: out <= 12'hb27;
      20'h03d2f: out <= 12'hb27;
      20'h03d30: out <= 12'hb27;
      20'h03d31: out <= 12'hb27;
      20'h03d32: out <= 12'hb27;
      20'h03d33: out <= 12'hb27;
      20'h03d34: out <= 12'hb27;
      20'h03d35: out <= 12'hb27;
      20'h03d36: out <= 12'hb27;
      20'h03d37: out <= 12'hb27;
      20'h03d38: out <= 12'hb27;
      20'h03d39: out <= 12'hb27;
      20'h03d3a: out <= 12'hb27;
      20'h03d3b: out <= 12'hb27;
      20'h03d3c: out <= 12'hb27;
      20'h03d3d: out <= 12'hb27;
      20'h03d3e: out <= 12'hb27;
      20'h03d3f: out <= 12'hb27;
      20'h03d40: out <= 12'hfff;
      20'h03d41: out <= 12'hc7f;
      20'h03d42: out <= 12'h72f;
      20'h03d43: out <= 12'hfff;
      20'h03d44: out <= 12'h72f;
      20'h03d45: out <= 12'hc7f;
      20'h03d46: out <= 12'hfff;
      20'h03d47: out <= 12'hfff;
      20'h03d48: out <= 12'hc7f;
      20'h03d49: out <= 12'h72f;
      20'h03d4a: out <= 12'h72f;
      20'h03d4b: out <= 12'hc7f;
      20'h03d4c: out <= 12'hfff;
      20'h03d4d: out <= 12'h72f;
      20'h03d4e: out <= 12'h72f;
      20'h03d4f: out <= 12'hc7f;
      20'h03d50: out <= 12'h72f;
      20'h03d51: out <= 12'hc7f;
      20'h03d52: out <= 12'hfff;
      20'h03d53: out <= 12'hfff;
      20'h03d54: out <= 12'h72f;
      20'h03d55: out <= 12'hc7f;
      20'h03d56: out <= 12'hfff;
      20'h03d57: out <= 12'hfff;
      20'h03d58: out <= 12'hc7f;
      20'h03d59: out <= 12'h72f;
      20'h03d5a: out <= 12'hfff;
      20'h03d5b: out <= 12'hc7f;
      20'h03d5c: out <= 12'h72f;
      20'h03d5d: out <= 12'h72f;
      20'h03d5e: out <= 12'h72f;
      20'h03d5f: out <= 12'hc7f;
      20'h03d60: out <= 12'h000;
      20'h03d61: out <= 12'hfff;
      20'h03d62: out <= 12'hc7f;
      20'h03d63: out <= 12'h72f;
      20'h03d64: out <= 12'h72f;
      20'h03d65: out <= 12'h72f;
      20'h03d66: out <= 12'hc7f;
      20'h03d67: out <= 12'hfff;
      20'h03d68: out <= 12'hfff;
      20'h03d69: out <= 12'hfff;
      20'h03d6a: out <= 12'hc7f;
      20'h03d6b: out <= 12'h72f;
      20'h03d6c: out <= 12'h72f;
      20'h03d6d: out <= 12'h72f;
      20'h03d6e: out <= 12'hc7f;
      20'h03d6f: out <= 12'hfff;
      20'h03d70: out <= 12'h222;
      20'h03d71: out <= 12'h72f;
      20'h03d72: out <= 12'hc7f;
      20'h03d73: out <= 12'hfff;
      20'h03d74: out <= 12'h72f;
      20'h03d75: out <= 12'h72f;
      20'h03d76: out <= 12'hc7f;
      20'h03d77: out <= 12'hfff;
      20'h03d78: out <= 12'hfff;
      20'h03d79: out <= 12'hfff;
      20'h03d7a: out <= 12'hc7f;
      20'h03d7b: out <= 12'h72f;
      20'h03d7c: out <= 12'h72f;
      20'h03d7d: out <= 12'hfff;
      20'h03d7e: out <= 12'hc7f;
      20'h03d7f: out <= 12'h72f;
      20'h03d80: out <= 12'hc7f;
      20'h03d81: out <= 12'h72f;
      20'h03d82: out <= 12'h72f;
      20'h03d83: out <= 12'hfff;
      20'h03d84: out <= 12'hc7f;
      20'h03d85: out <= 12'h72f;
      20'h03d86: out <= 12'h72f;
      20'h03d87: out <= 12'hc7f;
      20'h03d88: out <= 12'hfff;
      20'h03d89: out <= 12'hfff;
      20'h03d8a: out <= 12'hc7f;
      20'h03d8b: out <= 12'h72f;
      20'h03d8c: out <= 12'hfff;
      20'h03d8d: out <= 12'h72f;
      20'h03d8e: out <= 12'hc7f;
      20'h03d8f: out <= 12'hfff;
      20'h03d90: out <= 12'hc7f;
      20'h03d91: out <= 12'h72f;
      20'h03d92: out <= 12'h72f;
      20'h03d93: out <= 12'h72f;
      20'h03d94: out <= 12'hc7f;
      20'h03d95: out <= 12'hfff;
      20'h03d96: out <= 12'h72f;
      20'h03d97: out <= 12'hc7f;
      20'h03d98: out <= 12'hfff;
      20'h03d99: out <= 12'hfff;
      20'h03d9a: out <= 12'hc7f;
      20'h03d9b: out <= 12'h72f;
      20'h03d9c: out <= 12'hfff;
      20'h03d9d: out <= 12'hfff;
      20'h03d9e: out <= 12'hc7f;
      20'h03d9f: out <= 12'h72f;
      20'h03da0: out <= 12'h000;
      20'h03da1: out <= 12'hfff;
      20'h03da2: out <= 12'hc7f;
      20'h03da3: out <= 12'h72f;
      20'h03da4: out <= 12'h72f;
      20'h03da5: out <= 12'h72f;
      20'h03da6: out <= 12'h72f;
      20'h03da7: out <= 12'hc7f;
      20'h03da8: out <= 12'hfff;
      20'h03da9: out <= 12'hc7f;
      20'h03daa: out <= 12'h72f;
      20'h03dab: out <= 12'h72f;
      20'h03dac: out <= 12'h72f;
      20'h03dad: out <= 12'h72f;
      20'h03dae: out <= 12'hc7f;
      20'h03daf: out <= 12'hfff;
      20'h03db0: out <= 12'h222;
      20'h03db1: out <= 12'h72f;
      20'h03db2: out <= 12'hc7f;
      20'h03db3: out <= 12'hfff;
      20'h03db4: out <= 12'h72f;
      20'h03db5: out <= 12'h72f;
      20'h03db6: out <= 12'h72f;
      20'h03db7: out <= 12'hc7f;
      20'h03db8: out <= 12'hfff;
      20'h03db9: out <= 12'hc7f;
      20'h03dba: out <= 12'h72f;
      20'h03dbb: out <= 12'h72f;
      20'h03dbc: out <= 12'h72f;
      20'h03dbd: out <= 12'hfff;
      20'h03dbe: out <= 12'hc7f;
      20'h03dbf: out <= 12'h72f;
      20'h03dc0: out <= 12'h603;
      20'h03dc1: out <= 12'h603;
      20'h03dc2: out <= 12'h603;
      20'h03dc3: out <= 12'h603;
      20'h03dc4: out <= 12'h000;
      20'h03dc5: out <= 12'h000;
      20'h03dc6: out <= 12'hb27;
      20'h03dc7: out <= 12'hf87;
      20'h03dc8: out <= 12'hee9;
      20'h03dc9: out <= 12'hee9;
      20'h03dca: out <= 12'hee9;
      20'h03dcb: out <= 12'hee9;
      20'h03dcc: out <= 12'hee9;
      20'h03dcd: out <= 12'hee9;
      20'h03dce: out <= 12'hf87;
      20'h03dcf: out <= 12'hee9;
      20'h03dd0: out <= 12'hf87;
      20'h03dd1: out <= 12'hf87;
      20'h03dd2: out <= 12'hb27;
      20'h03dd3: out <= 12'h000;
      20'h03dd4: out <= 12'h000;
      20'h03dd5: out <= 12'hf87;
      20'h03dd6: out <= 12'hb27;
      20'h03dd7: out <= 12'hf87;
      20'h03dd8: out <= 12'hf87;
      20'h03dd9: out <= 12'hee9;
      20'h03dda: out <= 12'hf87;
      20'h03ddb: out <= 12'hf87;
      20'h03ddc: out <= 12'hf87;
      20'h03ddd: out <= 12'hb27;
      20'h03dde: out <= 12'hf87;
      20'h03ddf: out <= 12'hee9;
      20'h03de0: out <= 12'hf87;
      20'h03de1: out <= 12'hf87;
      20'h03de2: out <= 12'hee9;
      20'h03de3: out <= 12'hf87;
      20'h03de4: out <= 12'h000;
      20'h03de5: out <= 12'h000;
      20'h03de6: out <= 12'hb27;
      20'h03de7: out <= 12'hb27;
      20'h03de8: out <= 12'hb27;
      20'h03de9: out <= 12'hb27;
      20'h03dea: out <= 12'hf87;
      20'h03deb: out <= 12'hf87;
      20'h03dec: out <= 12'hf87;
      20'h03ded: out <= 12'hb27;
      20'h03dee: out <= 12'hf87;
      20'h03def: out <= 12'hee9;
      20'h03df0: out <= 12'hf87;
      20'h03df1: out <= 12'hb27;
      20'h03df2: out <= 12'hee9;
      20'h03df3: out <= 12'hf87;
      20'h03df4: out <= 12'h603;
      20'h03df5: out <= 12'h603;
      20'h03df6: out <= 12'h603;
      20'h03df7: out <= 12'h603;
      20'h03df8: out <= 12'h603;
      20'h03df9: out <= 12'h603;
      20'h03dfa: out <= 12'h603;
      20'h03dfb: out <= 12'h603;
      20'h03dfc: out <= 12'h603;
      20'h03dfd: out <= 12'h603;
      20'h03dfe: out <= 12'h603;
      20'h03dff: out <= 12'h603;
      20'h03e00: out <= 12'h603;
      20'h03e01: out <= 12'h603;
      20'h03e02: out <= 12'h603;
      20'h03e03: out <= 12'h603;
      20'h03e04: out <= 12'h603;
      20'h03e05: out <= 12'h603;
      20'h03e06: out <= 12'h603;
      20'h03e07: out <= 12'h603;
      20'h03e08: out <= 12'h603;
      20'h03e09: out <= 12'h603;
      20'h03e0a: out <= 12'h603;
      20'h03e0b: out <= 12'h603;
      20'h03e0c: out <= 12'h603;
      20'h03e0d: out <= 12'h603;
      20'h03e0e: out <= 12'h603;
      20'h03e0f: out <= 12'h603;
      20'h03e10: out <= 12'h603;
      20'h03e11: out <= 12'h603;
      20'h03e12: out <= 12'h603;
      20'h03e13: out <= 12'h603;
      20'h03e14: out <= 12'h603;
      20'h03e15: out <= 12'h603;
      20'h03e16: out <= 12'h603;
      20'h03e17: out <= 12'h603;
      20'h03e18: out <= 12'hee9;
      20'h03e19: out <= 12'hee9;
      20'h03e1a: out <= 12'hee9;
      20'h03e1b: out <= 12'hee9;
      20'h03e1c: out <= 12'hee9;
      20'h03e1d: out <= 12'hee9;
      20'h03e1e: out <= 12'hee9;
      20'h03e1f: out <= 12'hb27;
      20'h03e20: out <= 12'h000;
      20'h03e21: out <= 12'h000;
      20'h03e22: out <= 12'h000;
      20'h03e23: out <= 12'h000;
      20'h03e24: out <= 12'h000;
      20'h03e25: out <= 12'h000;
      20'h03e26: out <= 12'h000;
      20'h03e27: out <= 12'h000;
      20'h03e28: out <= 12'h000;
      20'h03e29: out <= 12'h000;
      20'h03e2a: out <= 12'h000;
      20'h03e2b: out <= 12'h000;
      20'h03e2c: out <= 12'h000;
      20'h03e2d: out <= 12'h000;
      20'h03e2e: out <= 12'h000;
      20'h03e2f: out <= 12'h000;
      20'h03e30: out <= 12'h000;
      20'h03e31: out <= 12'h000;
      20'h03e32: out <= 12'h000;
      20'h03e33: out <= 12'h000;
      20'h03e34: out <= 12'h000;
      20'h03e35: out <= 12'h000;
      20'h03e36: out <= 12'h000;
      20'h03e37: out <= 12'h000;
      20'h03e38: out <= 12'h000;
      20'h03e39: out <= 12'h000;
      20'h03e3a: out <= 12'h000;
      20'h03e3b: out <= 12'h000;
      20'h03e3c: out <= 12'h000;
      20'h03e3d: out <= 12'h000;
      20'h03e3e: out <= 12'h000;
      20'h03e3f: out <= 12'h000;
      20'h03e40: out <= 12'h000;
      20'h03e41: out <= 12'h000;
      20'h03e42: out <= 12'h000;
      20'h03e43: out <= 12'h000;
      20'h03e44: out <= 12'h000;
      20'h03e45: out <= 12'h000;
      20'h03e46: out <= 12'h000;
      20'h03e47: out <= 12'h000;
      20'h03e48: out <= 12'h000;
      20'h03e49: out <= 12'h000;
      20'h03e4a: out <= 12'h000;
      20'h03e4b: out <= 12'h000;
      20'h03e4c: out <= 12'h000;
      20'h03e4d: out <= 12'h000;
      20'h03e4e: out <= 12'h000;
      20'h03e4f: out <= 12'h000;
      20'h03e50: out <= 12'h000;
      20'h03e51: out <= 12'h000;
      20'h03e52: out <= 12'h000;
      20'h03e53: out <= 12'h000;
      20'h03e54: out <= 12'h000;
      20'h03e55: out <= 12'h000;
      20'h03e56: out <= 12'h000;
      20'h03e57: out <= 12'h000;
      20'h03e58: out <= 12'hfff;
      20'h03e59: out <= 12'hc7f;
      20'h03e5a: out <= 12'h72f;
      20'h03e5b: out <= 12'hc7f;
      20'h03e5c: out <= 12'h72f;
      20'h03e5d: out <= 12'h72f;
      20'h03e5e: out <= 12'hc7f;
      20'h03e5f: out <= 12'hc7f;
      20'h03e60: out <= 12'h72f;
      20'h03e61: out <= 12'h72f;
      20'h03e62: out <= 12'h72f;
      20'h03e63: out <= 12'hc7f;
      20'h03e64: out <= 12'hfff;
      20'h03e65: out <= 12'h000;
      20'h03e66: out <= 12'h000;
      20'h03e67: out <= 12'h000;
      20'h03e68: out <= 12'h72f;
      20'h03e69: out <= 12'hc7f;
      20'h03e6a: out <= 12'hfff;
      20'h03e6b: out <= 12'hc7f;
      20'h03e6c: out <= 12'h72f;
      20'h03e6d: out <= 12'h72f;
      20'h03e6e: out <= 12'hc7f;
      20'h03e6f: out <= 12'hc7f;
      20'h03e70: out <= 12'h72f;
      20'h03e71: out <= 12'h72f;
      20'h03e72: out <= 12'hfff;
      20'h03e73: out <= 12'hc7f;
      20'h03e74: out <= 12'h72f;
      20'h03e75: out <= 12'h222;
      20'h03e76: out <= 12'h222;
      20'h03e77: out <= 12'h222;
      20'h03e78: out <= 12'h000;
      20'h03e79: out <= 12'hfff;
      20'h03e7a: out <= 12'hc7f;
      20'h03e7b: out <= 12'h72f;
      20'h03e7c: out <= 12'h72f;
      20'h03e7d: out <= 12'h72f;
      20'h03e7e: out <= 12'hc7f;
      20'h03e7f: out <= 12'hfff;
      20'h03e80: out <= 12'hfff;
      20'h03e81: out <= 12'hfff;
      20'h03e82: out <= 12'hc7f;
      20'h03e83: out <= 12'h72f;
      20'h03e84: out <= 12'h72f;
      20'h03e85: out <= 12'h72f;
      20'h03e86: out <= 12'hc7f;
      20'h03e87: out <= 12'hfff;
      20'h03e88: out <= 12'h222;
      20'h03e89: out <= 12'h72f;
      20'h03e8a: out <= 12'hc7f;
      20'h03e8b: out <= 12'hfff;
      20'h03e8c: out <= 12'h72f;
      20'h03e8d: out <= 12'h72f;
      20'h03e8e: out <= 12'hc7f;
      20'h03e8f: out <= 12'hfff;
      20'h03e90: out <= 12'hfff;
      20'h03e91: out <= 12'hfff;
      20'h03e92: out <= 12'hc7f;
      20'h03e93: out <= 12'h72f;
      20'h03e94: out <= 12'h72f;
      20'h03e95: out <= 12'hfff;
      20'h03e96: out <= 12'hc7f;
      20'h03e97: out <= 12'h72f;
      20'h03e98: out <= 12'h000;
      20'h03e99: out <= 12'h000;
      20'h03e9a: out <= 12'h000;
      20'h03e9b: out <= 12'hfff;
      20'h03e9c: out <= 12'hc7f;
      20'h03e9d: out <= 12'h72f;
      20'h03e9e: out <= 12'h72f;
      20'h03e9f: out <= 12'h72f;
      20'h03ea0: out <= 12'hc7f;
      20'h03ea1: out <= 12'hc7f;
      20'h03ea2: out <= 12'h72f;
      20'h03ea3: out <= 12'h72f;
      20'h03ea4: out <= 12'hc7f;
      20'h03ea5: out <= 12'h72f;
      20'h03ea6: out <= 12'hc7f;
      20'h03ea7: out <= 12'hfff;
      20'h03ea8: out <= 12'h222;
      20'h03ea9: out <= 12'h222;
      20'h03eaa: out <= 12'h222;
      20'h03eab: out <= 12'h72f;
      20'h03eac: out <= 12'hc7f;
      20'h03ead: out <= 12'hfff;
      20'h03eae: out <= 12'h72f;
      20'h03eaf: out <= 12'h72f;
      20'h03eb0: out <= 12'hc7f;
      20'h03eb1: out <= 12'hc7f;
      20'h03eb2: out <= 12'h72f;
      20'h03eb3: out <= 12'h72f;
      20'h03eb4: out <= 12'hc7f;
      20'h03eb5: out <= 12'hfff;
      20'h03eb6: out <= 12'hc7f;
      20'h03eb7: out <= 12'h72f;
      20'h03eb8: out <= 12'h000;
      20'h03eb9: out <= 12'hc7f;
      20'h03eba: out <= 12'hfff;
      20'h03ebb: out <= 12'hc7f;
      20'h03ebc: out <= 12'h72f;
      20'h03ebd: out <= 12'h72f;
      20'h03ebe: out <= 12'h72f;
      20'h03ebf: out <= 12'h72f;
      20'h03ec0: out <= 12'h72f;
      20'h03ec1: out <= 12'h72f;
      20'h03ec2: out <= 12'h72f;
      20'h03ec3: out <= 12'h72f;
      20'h03ec4: out <= 12'h72f;
      20'h03ec5: out <= 12'hc7f;
      20'h03ec6: out <= 12'hfff;
      20'h03ec7: out <= 12'hc7f;
      20'h03ec8: out <= 12'h222;
      20'h03ec9: out <= 12'hc7f;
      20'h03eca: out <= 12'h72f;
      20'h03ecb: out <= 12'hc7f;
      20'h03ecc: out <= 12'hfff;
      20'h03ecd: out <= 12'hfff;
      20'h03ece: out <= 12'h72f;
      20'h03ecf: out <= 12'h72f;
      20'h03ed0: out <= 12'h72f;
      20'h03ed1: out <= 12'h72f;
      20'h03ed2: out <= 12'h72f;
      20'h03ed3: out <= 12'hfff;
      20'h03ed4: out <= 12'hfff;
      20'h03ed5: out <= 12'hc7f;
      20'h03ed6: out <= 12'h72f;
      20'h03ed7: out <= 12'hc7f;
      20'h03ed8: out <= 12'h603;
      20'h03ed9: out <= 12'h603;
      20'h03eda: out <= 12'h603;
      20'h03edb: out <= 12'h603;
      20'h03edc: out <= 12'h000;
      20'h03edd: out <= 12'h000;
      20'h03ede: out <= 12'hb27;
      20'h03edf: out <= 12'hf87;
      20'h03ee0: out <= 12'hee9;
      20'h03ee1: out <= 12'hee9;
      20'h03ee2: out <= 12'hee9;
      20'h03ee3: out <= 12'hee9;
      20'h03ee4: out <= 12'hee9;
      20'h03ee5: out <= 12'hf87;
      20'h03ee6: out <= 12'hee9;
      20'h03ee7: out <= 12'hf87;
      20'h03ee8: out <= 12'hf87;
      20'h03ee9: out <= 12'hb27;
      20'h03eea: out <= 12'hb27;
      20'h03eeb: out <= 12'h000;
      20'h03eec: out <= 12'h000;
      20'h03eed: out <= 12'hf87;
      20'h03eee: out <= 12'hb27;
      20'h03eef: out <= 12'hf87;
      20'h03ef0: out <= 12'hee9;
      20'h03ef1: out <= 12'hf87;
      20'h03ef2: out <= 12'hf87;
      20'h03ef3: out <= 12'hf87;
      20'h03ef4: out <= 12'hb27;
      20'h03ef5: out <= 12'hf87;
      20'h03ef6: out <= 12'hf87;
      20'h03ef7: out <= 12'hf87;
      20'h03ef8: out <= 12'hee9;
      20'h03ef9: out <= 12'hf87;
      20'h03efa: out <= 12'hee9;
      20'h03efb: out <= 12'hf87;
      20'h03efc: out <= 12'h000;
      20'h03efd: out <= 12'hf87;
      20'h03efe: out <= 12'hb27;
      20'h03eff: out <= 12'hb27;
      20'h03f00: out <= 12'hee9;
      20'h03f01: out <= 12'hf87;
      20'h03f02: out <= 12'hb27;
      20'h03f03: out <= 12'hb27;
      20'h03f04: out <= 12'hb27;
      20'h03f05: out <= 12'hf87;
      20'h03f06: out <= 12'hf87;
      20'h03f07: out <= 12'hf87;
      20'h03f08: out <= 12'hee9;
      20'h03f09: out <= 12'hf87;
      20'h03f0a: out <= 12'hee9;
      20'h03f0b: out <= 12'hf87;
      20'h03f0c: out <= 12'h603;
      20'h03f0d: out <= 12'h603;
      20'h03f0e: out <= 12'h603;
      20'h03f0f: out <= 12'h603;
      20'h03f10: out <= 12'h603;
      20'h03f11: out <= 12'h603;
      20'h03f12: out <= 12'h603;
      20'h03f13: out <= 12'h603;
      20'h03f14: out <= 12'h603;
      20'h03f15: out <= 12'h603;
      20'h03f16: out <= 12'h603;
      20'h03f17: out <= 12'h603;
      20'h03f18: out <= 12'h603;
      20'h03f19: out <= 12'h603;
      20'h03f1a: out <= 12'h603;
      20'h03f1b: out <= 12'h603;
      20'h03f1c: out <= 12'h603;
      20'h03f1d: out <= 12'h603;
      20'h03f1e: out <= 12'h603;
      20'h03f1f: out <= 12'h603;
      20'h03f20: out <= 12'h603;
      20'h03f21: out <= 12'h603;
      20'h03f22: out <= 12'h603;
      20'h03f23: out <= 12'h603;
      20'h03f24: out <= 12'h603;
      20'h03f25: out <= 12'h603;
      20'h03f26: out <= 12'h603;
      20'h03f27: out <= 12'h603;
      20'h03f28: out <= 12'h603;
      20'h03f29: out <= 12'h603;
      20'h03f2a: out <= 12'h603;
      20'h03f2b: out <= 12'h603;
      20'h03f2c: out <= 12'h603;
      20'h03f2d: out <= 12'h603;
      20'h03f2e: out <= 12'h603;
      20'h03f2f: out <= 12'h603;
      20'h03f30: out <= 12'hee9;
      20'h03f31: out <= 12'hf87;
      20'h03f32: out <= 12'hf87;
      20'h03f33: out <= 12'hf87;
      20'h03f34: out <= 12'hf87;
      20'h03f35: out <= 12'hf87;
      20'h03f36: out <= 12'hf87;
      20'h03f37: out <= 12'hb27;
      20'h03f38: out <= 12'h000;
      20'h03f39: out <= 12'h000;
      20'h03f3a: out <= 12'h000;
      20'h03f3b: out <= 12'h000;
      20'h03f3c: out <= 12'h000;
      20'h03f3d: out <= 12'h000;
      20'h03f3e: out <= 12'h000;
      20'h03f3f: out <= 12'h000;
      20'h03f40: out <= 12'h000;
      20'h03f41: out <= 12'h000;
      20'h03f42: out <= 12'h000;
      20'h03f43: out <= 12'h000;
      20'h03f44: out <= 12'h000;
      20'h03f45: out <= 12'h000;
      20'h03f46: out <= 12'h000;
      20'h03f47: out <= 12'h000;
      20'h03f48: out <= 12'h000;
      20'h03f49: out <= 12'h000;
      20'h03f4a: out <= 12'h000;
      20'h03f4b: out <= 12'h000;
      20'h03f4c: out <= 12'h000;
      20'h03f4d: out <= 12'h000;
      20'h03f4e: out <= 12'h000;
      20'h03f4f: out <= 12'h000;
      20'h03f50: out <= 12'h000;
      20'h03f51: out <= 12'h000;
      20'h03f52: out <= 12'h000;
      20'h03f53: out <= 12'h000;
      20'h03f54: out <= 12'h000;
      20'h03f55: out <= 12'h000;
      20'h03f56: out <= 12'h000;
      20'h03f57: out <= 12'h000;
      20'h03f58: out <= 12'h000;
      20'h03f59: out <= 12'h000;
      20'h03f5a: out <= 12'h000;
      20'h03f5b: out <= 12'h000;
      20'h03f5c: out <= 12'h000;
      20'h03f5d: out <= 12'h000;
      20'h03f5e: out <= 12'h000;
      20'h03f5f: out <= 12'h000;
      20'h03f60: out <= 12'h000;
      20'h03f61: out <= 12'h000;
      20'h03f62: out <= 12'h000;
      20'h03f63: out <= 12'h000;
      20'h03f64: out <= 12'h000;
      20'h03f65: out <= 12'h000;
      20'h03f66: out <= 12'h000;
      20'h03f67: out <= 12'h000;
      20'h03f68: out <= 12'h000;
      20'h03f69: out <= 12'h000;
      20'h03f6a: out <= 12'h000;
      20'h03f6b: out <= 12'h000;
      20'h03f6c: out <= 12'h000;
      20'h03f6d: out <= 12'h000;
      20'h03f6e: out <= 12'h000;
      20'h03f6f: out <= 12'h000;
      20'h03f70: out <= 12'h000;
      20'h03f71: out <= 12'hfff;
      20'h03f72: out <= 12'hc7f;
      20'h03f73: out <= 12'h72f;
      20'h03f74: out <= 12'hc7f;
      20'h03f75: out <= 12'h72f;
      20'h03f76: out <= 12'h72f;
      20'h03f77: out <= 12'h72f;
      20'h03f78: out <= 12'h72f;
      20'h03f79: out <= 12'h72f;
      20'h03f7a: out <= 12'hc7f;
      20'h03f7b: out <= 12'hfff;
      20'h03f7c: out <= 12'h000;
      20'h03f7d: out <= 12'h000;
      20'h03f7e: out <= 12'h000;
      20'h03f7f: out <= 12'h000;
      20'h03f80: out <= 12'h222;
      20'h03f81: out <= 12'h72f;
      20'h03f82: out <= 12'hc7f;
      20'h03f83: out <= 12'hfff;
      20'h03f84: out <= 12'hc7f;
      20'h03f85: out <= 12'h72f;
      20'h03f86: out <= 12'h72f;
      20'h03f87: out <= 12'h72f;
      20'h03f88: out <= 12'h72f;
      20'h03f89: out <= 12'hfff;
      20'h03f8a: out <= 12'hc7f;
      20'h03f8b: out <= 12'h72f;
      20'h03f8c: out <= 12'h222;
      20'h03f8d: out <= 12'h222;
      20'h03f8e: out <= 12'h222;
      20'h03f8f: out <= 12'h222;
      20'h03f90: out <= 12'h000;
      20'h03f91: out <= 12'hfff;
      20'h03f92: out <= 12'hc7f;
      20'h03f93: out <= 12'h72f;
      20'h03f94: out <= 12'h72f;
      20'h03f95: out <= 12'h72f;
      20'h03f96: out <= 12'h72f;
      20'h03f97: out <= 12'hc7f;
      20'h03f98: out <= 12'hfff;
      20'h03f99: out <= 12'hc7f;
      20'h03f9a: out <= 12'h72f;
      20'h03f9b: out <= 12'h72f;
      20'h03f9c: out <= 12'h72f;
      20'h03f9d: out <= 12'h72f;
      20'h03f9e: out <= 12'hc7f;
      20'h03f9f: out <= 12'hfff;
      20'h03fa0: out <= 12'h222;
      20'h03fa1: out <= 12'h72f;
      20'h03fa2: out <= 12'hc7f;
      20'h03fa3: out <= 12'hfff;
      20'h03fa4: out <= 12'h72f;
      20'h03fa5: out <= 12'h72f;
      20'h03fa6: out <= 12'h72f;
      20'h03fa7: out <= 12'hc7f;
      20'h03fa8: out <= 12'hfff;
      20'h03fa9: out <= 12'hc7f;
      20'h03faa: out <= 12'h72f;
      20'h03fab: out <= 12'h72f;
      20'h03fac: out <= 12'h72f;
      20'h03fad: out <= 12'hfff;
      20'h03fae: out <= 12'hc7f;
      20'h03faf: out <= 12'h72f;
      20'h03fb0: out <= 12'h000;
      20'h03fb1: out <= 12'h000;
      20'h03fb2: out <= 12'h000;
      20'h03fb3: out <= 12'h000;
      20'h03fb4: out <= 12'hfff;
      20'h03fb5: out <= 12'hc7f;
      20'h03fb6: out <= 12'h72f;
      20'h03fb7: out <= 12'h72f;
      20'h03fb8: out <= 12'h72f;
      20'h03fb9: out <= 12'h72f;
      20'h03fba: out <= 12'h72f;
      20'h03fbb: out <= 12'hc7f;
      20'h03fbc: out <= 12'h72f;
      20'h03fbd: out <= 12'hc7f;
      20'h03fbe: out <= 12'hfff;
      20'h03fbf: out <= 12'h000;
      20'h03fc0: out <= 12'h222;
      20'h03fc1: out <= 12'h222;
      20'h03fc2: out <= 12'h222;
      20'h03fc3: out <= 12'h222;
      20'h03fc4: out <= 12'h72f;
      20'h03fc5: out <= 12'hc7f;
      20'h03fc6: out <= 12'hfff;
      20'h03fc7: out <= 12'h72f;
      20'h03fc8: out <= 12'h72f;
      20'h03fc9: out <= 12'h72f;
      20'h03fca: out <= 12'h72f;
      20'h03fcb: out <= 12'hc7f;
      20'h03fcc: out <= 12'hfff;
      20'h03fcd: out <= 12'hc7f;
      20'h03fce: out <= 12'h72f;
      20'h03fcf: out <= 12'h222;
      20'h03fd0: out <= 12'h000;
      20'h03fd1: out <= 12'hc7f;
      20'h03fd2: out <= 12'h72f;
      20'h03fd3: out <= 12'hfff;
      20'h03fd4: out <= 12'hc7f;
      20'h03fd5: out <= 12'hc7f;
      20'h03fd6: out <= 12'h72f;
      20'h03fd7: out <= 12'h72f;
      20'h03fd8: out <= 12'h72f;
      20'h03fd9: out <= 12'h72f;
      20'h03fda: out <= 12'h72f;
      20'h03fdb: out <= 12'hc7f;
      20'h03fdc: out <= 12'hc7f;
      20'h03fdd: out <= 12'hfff;
      20'h03fde: out <= 12'h72f;
      20'h03fdf: out <= 12'hc7f;
      20'h03fe0: out <= 12'h222;
      20'h03fe1: out <= 12'hc7f;
      20'h03fe2: out <= 12'h72f;
      20'h03fe3: out <= 12'h72f;
      20'h03fe4: out <= 12'hc7f;
      20'h03fe5: out <= 12'hc7f;
      20'h03fe6: out <= 12'hfff;
      20'h03fe7: out <= 12'hfff;
      20'h03fe8: out <= 12'hfff;
      20'h03fe9: out <= 12'hfff;
      20'h03fea: out <= 12'hfff;
      20'h03feb: out <= 12'hc7f;
      20'h03fec: out <= 12'hc7f;
      20'h03fed: out <= 12'h72f;
      20'h03fee: out <= 12'h72f;
      20'h03fef: out <= 12'hc7f;
      20'h03ff0: out <= 12'h603;
      20'h03ff1: out <= 12'h603;
      20'h03ff2: out <= 12'h603;
      20'h03ff3: out <= 12'h603;
      20'h03ff4: out <= 12'h000;
      20'h03ff5: out <= 12'h000;
      20'h03ff6: out <= 12'hb27;
      20'h03ff7: out <= 12'hf87;
      20'h03ff8: out <= 12'hee9;
      20'h03ff9: out <= 12'hee9;
      20'h03ffa: out <= 12'hee9;
      20'h03ffb: out <= 12'hee9;
      20'h03ffc: out <= 12'hf87;
      20'h03ffd: out <= 12'hee9;
      20'h03ffe: out <= 12'hf87;
      20'h03fff: out <= 12'hf87;
      20'h04000: out <= 12'hb27;
      20'h04001: out <= 12'hf87;
      20'h04002: out <= 12'hb27;
      20'h04003: out <= 12'h000;
      20'h04004: out <= 12'h000;
      20'h04005: out <= 12'hf87;
      20'h04006: out <= 12'hb27;
      20'h04007: out <= 12'hee9;
      20'h04008: out <= 12'hf87;
      20'h04009: out <= 12'hf87;
      20'h0400a: out <= 12'hf87;
      20'h0400b: out <= 12'hb27;
      20'h0400c: out <= 12'hf87;
      20'h0400d: out <= 12'hb27;
      20'h0400e: out <= 12'hf87;
      20'h0400f: out <= 12'hf87;
      20'h04010: out <= 12'hf87;
      20'h04011: out <= 12'hee9;
      20'h04012: out <= 12'hee9;
      20'h04013: out <= 12'hf87;
      20'h04014: out <= 12'h000;
      20'h04015: out <= 12'hf87;
      20'h04016: out <= 12'hb27;
      20'h04017: out <= 12'hee9;
      20'h04018: out <= 12'hf87;
      20'h04019: out <= 12'hf87;
      20'h0401a: out <= 12'hf87;
      20'h0401b: out <= 12'hb27;
      20'h0401c: out <= 12'hf87;
      20'h0401d: out <= 12'hb27;
      20'h0401e: out <= 12'hf87;
      20'h0401f: out <= 12'hf87;
      20'h04020: out <= 12'hf87;
      20'h04021: out <= 12'hee9;
      20'h04022: out <= 12'hee9;
      20'h04023: out <= 12'hf87;
      20'h04024: out <= 12'h603;
      20'h04025: out <= 12'h603;
      20'h04026: out <= 12'h603;
      20'h04027: out <= 12'h603;
      20'h04028: out <= 12'h603;
      20'h04029: out <= 12'h603;
      20'h0402a: out <= 12'h603;
      20'h0402b: out <= 12'h603;
      20'h0402c: out <= 12'h603;
      20'h0402d: out <= 12'h603;
      20'h0402e: out <= 12'h603;
      20'h0402f: out <= 12'h603;
      20'h04030: out <= 12'h603;
      20'h04031: out <= 12'h603;
      20'h04032: out <= 12'h603;
      20'h04033: out <= 12'h603;
      20'h04034: out <= 12'h603;
      20'h04035: out <= 12'h603;
      20'h04036: out <= 12'h603;
      20'h04037: out <= 12'h603;
      20'h04038: out <= 12'h603;
      20'h04039: out <= 12'h603;
      20'h0403a: out <= 12'h603;
      20'h0403b: out <= 12'h603;
      20'h0403c: out <= 12'h603;
      20'h0403d: out <= 12'h603;
      20'h0403e: out <= 12'h603;
      20'h0403f: out <= 12'h603;
      20'h04040: out <= 12'h603;
      20'h04041: out <= 12'h603;
      20'h04042: out <= 12'h603;
      20'h04043: out <= 12'h603;
      20'h04044: out <= 12'h603;
      20'h04045: out <= 12'h603;
      20'h04046: out <= 12'h603;
      20'h04047: out <= 12'h603;
      20'h04048: out <= 12'hee9;
      20'h04049: out <= 12'hf87;
      20'h0404a: out <= 12'hee9;
      20'h0404b: out <= 12'hee9;
      20'h0404c: out <= 12'hee9;
      20'h0404d: out <= 12'hb27;
      20'h0404e: out <= 12'hf87;
      20'h0404f: out <= 12'hb27;
      20'h04050: out <= 12'h000;
      20'h04051: out <= 12'h000;
      20'h04052: out <= 12'h000;
      20'h04053: out <= 12'h000;
      20'h04054: out <= 12'h000;
      20'h04055: out <= 12'h000;
      20'h04056: out <= 12'h000;
      20'h04057: out <= 12'h000;
      20'h04058: out <= 12'h000;
      20'h04059: out <= 12'h000;
      20'h0405a: out <= 12'h000;
      20'h0405b: out <= 12'h000;
      20'h0405c: out <= 12'h000;
      20'h0405d: out <= 12'h000;
      20'h0405e: out <= 12'h000;
      20'h0405f: out <= 12'h000;
      20'h04060: out <= 12'h000;
      20'h04061: out <= 12'h000;
      20'h04062: out <= 12'h000;
      20'h04063: out <= 12'h000;
      20'h04064: out <= 12'h000;
      20'h04065: out <= 12'h000;
      20'h04066: out <= 12'h000;
      20'h04067: out <= 12'h000;
      20'h04068: out <= 12'h000;
      20'h04069: out <= 12'h000;
      20'h0406a: out <= 12'h000;
      20'h0406b: out <= 12'h000;
      20'h0406c: out <= 12'h000;
      20'h0406d: out <= 12'h000;
      20'h0406e: out <= 12'h000;
      20'h0406f: out <= 12'h000;
      20'h04070: out <= 12'h000;
      20'h04071: out <= 12'h000;
      20'h04072: out <= 12'h000;
      20'h04073: out <= 12'h000;
      20'h04074: out <= 12'h000;
      20'h04075: out <= 12'h000;
      20'h04076: out <= 12'h000;
      20'h04077: out <= 12'h000;
      20'h04078: out <= 12'h000;
      20'h04079: out <= 12'h000;
      20'h0407a: out <= 12'h000;
      20'h0407b: out <= 12'h000;
      20'h0407c: out <= 12'h000;
      20'h0407d: out <= 12'h000;
      20'h0407e: out <= 12'h000;
      20'h0407f: out <= 12'h000;
      20'h04080: out <= 12'h000;
      20'h04081: out <= 12'h000;
      20'h04082: out <= 12'h000;
      20'h04083: out <= 12'h000;
      20'h04084: out <= 12'h000;
      20'h04085: out <= 12'h000;
      20'h04086: out <= 12'h000;
      20'h04087: out <= 12'h000;
      20'h04088: out <= 12'h000;
      20'h04089: out <= 12'hfff;
      20'h0408a: out <= 12'hc7f;
      20'h0408b: out <= 12'h72f;
      20'h0408c: out <= 12'h72f;
      20'h0408d: out <= 12'h72f;
      20'h0408e: out <= 12'h72f;
      20'h0408f: out <= 12'h72f;
      20'h04090: out <= 12'h72f;
      20'h04091: out <= 12'h72f;
      20'h04092: out <= 12'hc7f;
      20'h04093: out <= 12'hfff;
      20'h04094: out <= 12'h000;
      20'h04095: out <= 12'h000;
      20'h04096: out <= 12'h000;
      20'h04097: out <= 12'h000;
      20'h04098: out <= 12'h222;
      20'h04099: out <= 12'h72f;
      20'h0409a: out <= 12'hc7f;
      20'h0409b: out <= 12'hfff;
      20'h0409c: out <= 12'h72f;
      20'h0409d: out <= 12'h72f;
      20'h0409e: out <= 12'h72f;
      20'h0409f: out <= 12'h72f;
      20'h040a0: out <= 12'h72f;
      20'h040a1: out <= 12'hfff;
      20'h040a2: out <= 12'hc7f;
      20'h040a3: out <= 12'h72f;
      20'h040a4: out <= 12'h222;
      20'h040a5: out <= 12'h222;
      20'h040a6: out <= 12'h222;
      20'h040a7: out <= 12'h222;
      20'h040a8: out <= 12'h000;
      20'h040a9: out <= 12'hfff;
      20'h040aa: out <= 12'hc7f;
      20'h040ab: out <= 12'h72f;
      20'h040ac: out <= 12'h72f;
      20'h040ad: out <= 12'hc7f;
      20'h040ae: out <= 12'h72f;
      20'h040af: out <= 12'h72f;
      20'h040b0: out <= 12'h72f;
      20'h040b1: out <= 12'h72f;
      20'h040b2: out <= 12'h72f;
      20'h040b3: out <= 12'hc7f;
      20'h040b4: out <= 12'h72f;
      20'h040b5: out <= 12'h72f;
      20'h040b6: out <= 12'hc7f;
      20'h040b7: out <= 12'hfff;
      20'h040b8: out <= 12'h222;
      20'h040b9: out <= 12'h72f;
      20'h040ba: out <= 12'hc7f;
      20'h040bb: out <= 12'hfff;
      20'h040bc: out <= 12'h72f;
      20'h040bd: out <= 12'hc7f;
      20'h040be: out <= 12'h72f;
      20'h040bf: out <= 12'h72f;
      20'h040c0: out <= 12'h72f;
      20'h040c1: out <= 12'h72f;
      20'h040c2: out <= 12'h72f;
      20'h040c3: out <= 12'hc7f;
      20'h040c4: out <= 12'h72f;
      20'h040c5: out <= 12'hfff;
      20'h040c6: out <= 12'hc7f;
      20'h040c7: out <= 12'h72f;
      20'h040c8: out <= 12'h000;
      20'h040c9: out <= 12'h000;
      20'h040ca: out <= 12'h000;
      20'h040cb: out <= 12'h000;
      20'h040cc: out <= 12'hfff;
      20'h040cd: out <= 12'hc7f;
      20'h040ce: out <= 12'h72f;
      20'h040cf: out <= 12'h72f;
      20'h040d0: out <= 12'h72f;
      20'h040d1: out <= 12'h72f;
      20'h040d2: out <= 12'h72f;
      20'h040d3: out <= 12'h72f;
      20'h040d4: out <= 12'h72f;
      20'h040d5: out <= 12'hc7f;
      20'h040d6: out <= 12'hfff;
      20'h040d7: out <= 12'h000;
      20'h040d8: out <= 12'h222;
      20'h040d9: out <= 12'h222;
      20'h040da: out <= 12'h222;
      20'h040db: out <= 12'h222;
      20'h040dc: out <= 12'h72f;
      20'h040dd: out <= 12'hc7f;
      20'h040de: out <= 12'hfff;
      20'h040df: out <= 12'h72f;
      20'h040e0: out <= 12'h72f;
      20'h040e1: out <= 12'h72f;
      20'h040e2: out <= 12'h72f;
      20'h040e3: out <= 12'h72f;
      20'h040e4: out <= 12'hfff;
      20'h040e5: out <= 12'hc7f;
      20'h040e6: out <= 12'h72f;
      20'h040e7: out <= 12'h222;
      20'h040e8: out <= 12'h000;
      20'h040e9: out <= 12'hfff;
      20'h040ea: out <= 12'hfff;
      20'h040eb: out <= 12'hfff;
      20'h040ec: out <= 12'hfff;
      20'h040ed: out <= 12'hfff;
      20'h040ee: out <= 12'hc7f;
      20'h040ef: out <= 12'hc7f;
      20'h040f0: out <= 12'hc7f;
      20'h040f1: out <= 12'hc7f;
      20'h040f2: out <= 12'hc7f;
      20'h040f3: out <= 12'hfff;
      20'h040f4: out <= 12'hfff;
      20'h040f5: out <= 12'hfff;
      20'h040f6: out <= 12'hfff;
      20'h040f7: out <= 12'hfff;
      20'h040f8: out <= 12'h222;
      20'h040f9: out <= 12'hfff;
      20'h040fa: out <= 12'hfff;
      20'h040fb: out <= 12'hfff;
      20'h040fc: out <= 12'h72f;
      20'h040fd: out <= 12'h72f;
      20'h040fe: out <= 12'hc7f;
      20'h040ff: out <= 12'hc7f;
      20'h04100: out <= 12'hc7f;
      20'h04101: out <= 12'hc7f;
      20'h04102: out <= 12'hc7f;
      20'h04103: out <= 12'h72f;
      20'h04104: out <= 12'h72f;
      20'h04105: out <= 12'hfff;
      20'h04106: out <= 12'hfff;
      20'h04107: out <= 12'hfff;
      20'h04108: out <= 12'h603;
      20'h04109: out <= 12'h603;
      20'h0410a: out <= 12'h603;
      20'h0410b: out <= 12'h603;
      20'h0410c: out <= 12'h000;
      20'h0410d: out <= 12'h000;
      20'h0410e: out <= 12'hb27;
      20'h0410f: out <= 12'hf87;
      20'h04110: out <= 12'hf87;
      20'h04111: out <= 12'hee9;
      20'h04112: out <= 12'hee9;
      20'h04113: out <= 12'hf87;
      20'h04114: out <= 12'hee9;
      20'h04115: out <= 12'hf87;
      20'h04116: out <= 12'hf87;
      20'h04117: out <= 12'hb27;
      20'h04118: out <= 12'hf87;
      20'h04119: out <= 12'hb27;
      20'h0411a: out <= 12'hb27;
      20'h0411b: out <= 12'h000;
      20'h0411c: out <= 12'h000;
      20'h0411d: out <= 12'hf87;
      20'h0411e: out <= 12'hee9;
      20'h0411f: out <= 12'hf87;
      20'h04120: out <= 12'hf87;
      20'h04121: out <= 12'hf87;
      20'h04122: out <= 12'hb27;
      20'h04123: out <= 12'hf87;
      20'h04124: out <= 12'hf87;
      20'h04125: out <= 12'hf87;
      20'h04126: out <= 12'hb27;
      20'h04127: out <= 12'hf87;
      20'h04128: out <= 12'hf87;
      20'h04129: out <= 12'hf87;
      20'h0412a: out <= 12'hee9;
      20'h0412b: out <= 12'hf87;
      20'h0412c: out <= 12'h000;
      20'h0412d: out <= 12'hf87;
      20'h0412e: out <= 12'hee9;
      20'h0412f: out <= 12'hf87;
      20'h04130: out <= 12'hf87;
      20'h04131: out <= 12'hf87;
      20'h04132: out <= 12'hb27;
      20'h04133: out <= 12'hb27;
      20'h04134: out <= 12'hf87;
      20'h04135: out <= 12'hf87;
      20'h04136: out <= 12'hb27;
      20'h04137: out <= 12'hf87;
      20'h04138: out <= 12'hf87;
      20'h04139: out <= 12'hf87;
      20'h0413a: out <= 12'hee9;
      20'h0413b: out <= 12'hf87;
      20'h0413c: out <= 12'h603;
      20'h0413d: out <= 12'h603;
      20'h0413e: out <= 12'h603;
      20'h0413f: out <= 12'h603;
      20'h04140: out <= 12'h603;
      20'h04141: out <= 12'h603;
      20'h04142: out <= 12'h603;
      20'h04143: out <= 12'h603;
      20'h04144: out <= 12'h603;
      20'h04145: out <= 12'h603;
      20'h04146: out <= 12'h603;
      20'h04147: out <= 12'h603;
      20'h04148: out <= 12'h603;
      20'h04149: out <= 12'h603;
      20'h0414a: out <= 12'h603;
      20'h0414b: out <= 12'h603;
      20'h0414c: out <= 12'h603;
      20'h0414d: out <= 12'h603;
      20'h0414e: out <= 12'h603;
      20'h0414f: out <= 12'h603;
      20'h04150: out <= 12'h603;
      20'h04151: out <= 12'h603;
      20'h04152: out <= 12'h603;
      20'h04153: out <= 12'h603;
      20'h04154: out <= 12'h603;
      20'h04155: out <= 12'h603;
      20'h04156: out <= 12'h603;
      20'h04157: out <= 12'h603;
      20'h04158: out <= 12'h603;
      20'h04159: out <= 12'h603;
      20'h0415a: out <= 12'h603;
      20'h0415b: out <= 12'h603;
      20'h0415c: out <= 12'h603;
      20'h0415d: out <= 12'h603;
      20'h0415e: out <= 12'h603;
      20'h0415f: out <= 12'h603;
      20'h04160: out <= 12'hee9;
      20'h04161: out <= 12'hf87;
      20'h04162: out <= 12'hee9;
      20'h04163: out <= 12'hf87;
      20'h04164: out <= 12'hf87;
      20'h04165: out <= 12'hb27;
      20'h04166: out <= 12'hf87;
      20'h04167: out <= 12'hb27;
      20'h04168: out <= 12'h000;
      20'h04169: out <= 12'h000;
      20'h0416a: out <= 12'h000;
      20'h0416b: out <= 12'h000;
      20'h0416c: out <= 12'h000;
      20'h0416d: out <= 12'h000;
      20'h0416e: out <= 12'h000;
      20'h0416f: out <= 12'h000;
      20'h04170: out <= 12'h000;
      20'h04171: out <= 12'h000;
      20'h04172: out <= 12'h000;
      20'h04173: out <= 12'h000;
      20'h04174: out <= 12'h000;
      20'h04175: out <= 12'h000;
      20'h04176: out <= 12'h000;
      20'h04177: out <= 12'h000;
      20'h04178: out <= 12'h000;
      20'h04179: out <= 12'h000;
      20'h0417a: out <= 12'h000;
      20'h0417b: out <= 12'h000;
      20'h0417c: out <= 12'h000;
      20'h0417d: out <= 12'h000;
      20'h0417e: out <= 12'h000;
      20'h0417f: out <= 12'h000;
      20'h04180: out <= 12'h000;
      20'h04181: out <= 12'h000;
      20'h04182: out <= 12'h000;
      20'h04183: out <= 12'h000;
      20'h04184: out <= 12'h000;
      20'h04185: out <= 12'h000;
      20'h04186: out <= 12'h000;
      20'h04187: out <= 12'h000;
      20'h04188: out <= 12'h000;
      20'h04189: out <= 12'h000;
      20'h0418a: out <= 12'h000;
      20'h0418b: out <= 12'h000;
      20'h0418c: out <= 12'h000;
      20'h0418d: out <= 12'h000;
      20'h0418e: out <= 12'h000;
      20'h0418f: out <= 12'h000;
      20'h04190: out <= 12'h000;
      20'h04191: out <= 12'h000;
      20'h04192: out <= 12'h000;
      20'h04193: out <= 12'h000;
      20'h04194: out <= 12'h000;
      20'h04195: out <= 12'h000;
      20'h04196: out <= 12'h000;
      20'h04197: out <= 12'h000;
      20'h04198: out <= 12'h000;
      20'h04199: out <= 12'h000;
      20'h0419a: out <= 12'h000;
      20'h0419b: out <= 12'h000;
      20'h0419c: out <= 12'h000;
      20'h0419d: out <= 12'h000;
      20'h0419e: out <= 12'h000;
      20'h0419f: out <= 12'h000;
      20'h041a0: out <= 12'h000;
      20'h041a1: out <= 12'hc7f;
      20'h041a2: out <= 12'hfff;
      20'h041a3: out <= 12'hc7f;
      20'h041a4: out <= 12'h72f;
      20'h041a5: out <= 12'h72f;
      20'h041a6: out <= 12'h72f;
      20'h041a7: out <= 12'h72f;
      20'h041a8: out <= 12'h72f;
      20'h041a9: out <= 12'hc7f;
      20'h041aa: out <= 12'hfff;
      20'h041ab: out <= 12'hfff;
      20'h041ac: out <= 12'hc7f;
      20'h041ad: out <= 12'h000;
      20'h041ae: out <= 12'h000;
      20'h041af: out <= 12'h000;
      20'h041b0: out <= 12'h222;
      20'h041b1: out <= 12'hc7f;
      20'h041b2: out <= 12'hfff;
      20'h041b3: out <= 12'hc7f;
      20'h041b4: out <= 12'hfff;
      20'h041b5: out <= 12'hfff;
      20'h041b6: out <= 12'hfff;
      20'h041b7: out <= 12'hfff;
      20'h041b8: out <= 12'hfff;
      20'h041b9: out <= 12'hc7f;
      20'h041ba: out <= 12'h72f;
      20'h041bb: out <= 12'hfff;
      20'h041bc: out <= 12'hc7f;
      20'h041bd: out <= 12'h222;
      20'h041be: out <= 12'h222;
      20'h041bf: out <= 12'h222;
      20'h041c0: out <= 12'h000;
      20'h041c1: out <= 12'hc7f;
      20'h041c2: out <= 12'hfff;
      20'h041c3: out <= 12'hc7f;
      20'h041c4: out <= 12'h72f;
      20'h041c5: out <= 12'h72f;
      20'h041c6: out <= 12'hc7f;
      20'h041c7: out <= 12'hfff;
      20'h041c8: out <= 12'hfff;
      20'h041c9: out <= 12'hfff;
      20'h041ca: out <= 12'hc7f;
      20'h041cb: out <= 12'h72f;
      20'h041cc: out <= 12'h72f;
      20'h041cd: out <= 12'hc7f;
      20'h041ce: out <= 12'hfff;
      20'h041cf: out <= 12'hc7f;
      20'h041d0: out <= 12'h222;
      20'h041d1: out <= 12'hc7f;
      20'h041d2: out <= 12'h72f;
      20'h041d3: out <= 12'hc7f;
      20'h041d4: out <= 12'hfff;
      20'h041d5: out <= 12'hfff;
      20'h041d6: out <= 12'hc7f;
      20'h041d7: out <= 12'hfff;
      20'h041d8: out <= 12'hfff;
      20'h041d9: out <= 12'hfff;
      20'h041da: out <= 12'hc7f;
      20'h041db: out <= 12'hfff;
      20'h041dc: out <= 12'hfff;
      20'h041dd: out <= 12'hc7f;
      20'h041de: out <= 12'h72f;
      20'h041df: out <= 12'hc7f;
      20'h041e0: out <= 12'h000;
      20'h041e1: out <= 12'h000;
      20'h041e2: out <= 12'h000;
      20'h041e3: out <= 12'hc7f;
      20'h041e4: out <= 12'hfff;
      20'h041e5: out <= 12'hfff;
      20'h041e6: out <= 12'hc7f;
      20'h041e7: out <= 12'h72f;
      20'h041e8: out <= 12'h72f;
      20'h041e9: out <= 12'h72f;
      20'h041ea: out <= 12'h72f;
      20'h041eb: out <= 12'h72f;
      20'h041ec: out <= 12'hc7f;
      20'h041ed: out <= 12'hfff;
      20'h041ee: out <= 12'hc7f;
      20'h041ef: out <= 12'h000;
      20'h041f0: out <= 12'h222;
      20'h041f1: out <= 12'h222;
      20'h041f2: out <= 12'h222;
      20'h041f3: out <= 12'hc7f;
      20'h041f4: out <= 12'hfff;
      20'h041f5: out <= 12'h72f;
      20'h041f6: out <= 12'hc7f;
      20'h041f7: out <= 12'hfff;
      20'h041f8: out <= 12'hfff;
      20'h041f9: out <= 12'hfff;
      20'h041fa: out <= 12'hfff;
      20'h041fb: out <= 12'hfff;
      20'h041fc: out <= 12'hc7f;
      20'h041fd: out <= 12'hfff;
      20'h041fe: out <= 12'hc7f;
      20'h041ff: out <= 12'h222;
      20'h04200: out <= 12'h000;
      20'h04201: out <= 12'hc7f;
      20'h04202: out <= 12'h72f;
      20'h04203: out <= 12'hc7f;
      20'h04204: out <= 12'h000;
      20'h04205: out <= 12'h000;
      20'h04206: out <= 12'hfff;
      20'h04207: out <= 12'hfff;
      20'h04208: out <= 12'hfff;
      20'h04209: out <= 12'hfff;
      20'h0420a: out <= 12'hfff;
      20'h0420b: out <= 12'h000;
      20'h0420c: out <= 12'h000;
      20'h0420d: out <= 12'hc7f;
      20'h0420e: out <= 12'h72f;
      20'h0420f: out <= 12'hc7f;
      20'h04210: out <= 12'h222;
      20'h04211: out <= 12'hc7f;
      20'h04212: out <= 12'h72f;
      20'h04213: out <= 12'hc7f;
      20'h04214: out <= 12'h222;
      20'h04215: out <= 12'h222;
      20'h04216: out <= 12'h72f;
      20'h04217: out <= 12'h72f;
      20'h04218: out <= 12'h72f;
      20'h04219: out <= 12'h72f;
      20'h0421a: out <= 12'h72f;
      20'h0421b: out <= 12'h222;
      20'h0421c: out <= 12'h222;
      20'h0421d: out <= 12'hc7f;
      20'h0421e: out <= 12'h72f;
      20'h0421f: out <= 12'hc7f;
      20'h04220: out <= 12'h603;
      20'h04221: out <= 12'h603;
      20'h04222: out <= 12'h603;
      20'h04223: out <= 12'h603;
      20'h04224: out <= 12'h000;
      20'h04225: out <= 12'h000;
      20'h04226: out <= 12'hb27;
      20'h04227: out <= 12'hb27;
      20'h04228: out <= 12'hf87;
      20'h04229: out <= 12'hf87;
      20'h0422a: out <= 12'hf87;
      20'h0422b: out <= 12'hf87;
      20'h0422c: out <= 12'hf87;
      20'h0422d: out <= 12'hf87;
      20'h0422e: out <= 12'hb27;
      20'h0422f: out <= 12'hf87;
      20'h04230: out <= 12'hb27;
      20'h04231: out <= 12'hb27;
      20'h04232: out <= 12'hb27;
      20'h04233: out <= 12'h000;
      20'h04234: out <= 12'h000;
      20'h04235: out <= 12'hee9;
      20'h04236: out <= 12'hf87;
      20'h04237: out <= 12'hb27;
      20'h04238: out <= 12'hf87;
      20'h04239: out <= 12'hb27;
      20'h0423a: out <= 12'hf87;
      20'h0423b: out <= 12'hf87;
      20'h0423c: out <= 12'hf87;
      20'h0423d: out <= 12'hf87;
      20'h0423e: out <= 12'hf87;
      20'h0423f: out <= 12'hb27;
      20'h04240: out <= 12'hf87;
      20'h04241: out <= 12'hb27;
      20'h04242: out <= 12'hf87;
      20'h04243: out <= 12'hb27;
      20'h04244: out <= 12'h000;
      20'h04245: out <= 12'hee9;
      20'h04246: out <= 12'hf87;
      20'h04247: out <= 12'hb27;
      20'h04248: out <= 12'hf87;
      20'h04249: out <= 12'hb27;
      20'h0424a: out <= 12'hb27;
      20'h0424b: out <= 12'hb27;
      20'h0424c: out <= 12'hb27;
      20'h0424d: out <= 12'hf87;
      20'h0424e: out <= 12'hf87;
      20'h0424f: out <= 12'hb27;
      20'h04250: out <= 12'hf87;
      20'h04251: out <= 12'hb27;
      20'h04252: out <= 12'hf87;
      20'h04253: out <= 12'hb27;
      20'h04254: out <= 12'h603;
      20'h04255: out <= 12'h603;
      20'h04256: out <= 12'h603;
      20'h04257: out <= 12'h603;
      20'h04258: out <= 12'h603;
      20'h04259: out <= 12'h603;
      20'h0425a: out <= 12'h603;
      20'h0425b: out <= 12'h603;
      20'h0425c: out <= 12'h603;
      20'h0425d: out <= 12'h603;
      20'h0425e: out <= 12'h603;
      20'h0425f: out <= 12'h603;
      20'h04260: out <= 12'h603;
      20'h04261: out <= 12'h603;
      20'h04262: out <= 12'h603;
      20'h04263: out <= 12'h603;
      20'h04264: out <= 12'h603;
      20'h04265: out <= 12'h603;
      20'h04266: out <= 12'h603;
      20'h04267: out <= 12'h603;
      20'h04268: out <= 12'h603;
      20'h04269: out <= 12'h603;
      20'h0426a: out <= 12'h603;
      20'h0426b: out <= 12'h603;
      20'h0426c: out <= 12'h603;
      20'h0426d: out <= 12'h603;
      20'h0426e: out <= 12'h603;
      20'h0426f: out <= 12'h603;
      20'h04270: out <= 12'h603;
      20'h04271: out <= 12'h603;
      20'h04272: out <= 12'h603;
      20'h04273: out <= 12'h603;
      20'h04274: out <= 12'h603;
      20'h04275: out <= 12'h603;
      20'h04276: out <= 12'h603;
      20'h04277: out <= 12'h603;
      20'h04278: out <= 12'hee9;
      20'h04279: out <= 12'hf87;
      20'h0427a: out <= 12'hee9;
      20'h0427b: out <= 12'hf87;
      20'h0427c: out <= 12'hf87;
      20'h0427d: out <= 12'hb27;
      20'h0427e: out <= 12'hf87;
      20'h0427f: out <= 12'hb27;
      20'h04280: out <= 12'h000;
      20'h04281: out <= 12'h000;
      20'h04282: out <= 12'h000;
      20'h04283: out <= 12'h000;
      20'h04284: out <= 12'h000;
      20'h04285: out <= 12'h000;
      20'h04286: out <= 12'h000;
      20'h04287: out <= 12'h000;
      20'h04288: out <= 12'h000;
      20'h04289: out <= 12'h000;
      20'h0428a: out <= 12'h000;
      20'h0428b: out <= 12'h000;
      20'h0428c: out <= 12'h000;
      20'h0428d: out <= 12'h000;
      20'h0428e: out <= 12'h000;
      20'h0428f: out <= 12'h000;
      20'h04290: out <= 12'h000;
      20'h04291: out <= 12'h000;
      20'h04292: out <= 12'h000;
      20'h04293: out <= 12'h000;
      20'h04294: out <= 12'h000;
      20'h04295: out <= 12'h000;
      20'h04296: out <= 12'h000;
      20'h04297: out <= 12'h000;
      20'h04298: out <= 12'h000;
      20'h04299: out <= 12'h000;
      20'h0429a: out <= 12'h000;
      20'h0429b: out <= 12'h000;
      20'h0429c: out <= 12'h000;
      20'h0429d: out <= 12'h000;
      20'h0429e: out <= 12'h000;
      20'h0429f: out <= 12'h000;
      20'h042a0: out <= 12'h000;
      20'h042a1: out <= 12'h000;
      20'h042a2: out <= 12'h000;
      20'h042a3: out <= 12'h000;
      20'h042a4: out <= 12'h000;
      20'h042a5: out <= 12'h000;
      20'h042a6: out <= 12'h000;
      20'h042a7: out <= 12'h000;
      20'h042a8: out <= 12'h000;
      20'h042a9: out <= 12'h000;
      20'h042aa: out <= 12'h000;
      20'h042ab: out <= 12'h000;
      20'h042ac: out <= 12'h000;
      20'h042ad: out <= 12'h000;
      20'h042ae: out <= 12'h000;
      20'h042af: out <= 12'h000;
      20'h042b0: out <= 12'h000;
      20'h042b1: out <= 12'h000;
      20'h042b2: out <= 12'h000;
      20'h042b3: out <= 12'h000;
      20'h042b4: out <= 12'h000;
      20'h042b5: out <= 12'h000;
      20'h042b6: out <= 12'h000;
      20'h042b7: out <= 12'h000;
      20'h042b8: out <= 12'h000;
      20'h042b9: out <= 12'h72f;
      20'h042ba: out <= 12'hfff;
      20'h042bb: out <= 12'hfff;
      20'h042bc: out <= 12'hc7f;
      20'h042bd: out <= 12'hc7f;
      20'h042be: out <= 12'hc7f;
      20'h042bf: out <= 12'hc7f;
      20'h042c0: out <= 12'hc7f;
      20'h042c1: out <= 12'hfff;
      20'h042c2: out <= 12'h72f;
      20'h042c3: out <= 12'hfff;
      20'h042c4: out <= 12'h72f;
      20'h042c5: out <= 12'h000;
      20'h042c6: out <= 12'h000;
      20'h042c7: out <= 12'h000;
      20'h042c8: out <= 12'h222;
      20'h042c9: out <= 12'h72f;
      20'h042ca: out <= 12'hfff;
      20'h042cb: out <= 12'h72f;
      20'h042cc: out <= 12'hc7f;
      20'h042cd: out <= 12'hc7f;
      20'h042ce: out <= 12'hc7f;
      20'h042cf: out <= 12'hc7f;
      20'h042d0: out <= 12'hc7f;
      20'h042d1: out <= 12'h72f;
      20'h042d2: out <= 12'h72f;
      20'h042d3: out <= 12'hfff;
      20'h042d4: out <= 12'h72f;
      20'h042d5: out <= 12'h222;
      20'h042d6: out <= 12'h222;
      20'h042d7: out <= 12'h222;
      20'h042d8: out <= 12'h000;
      20'h042d9: out <= 12'hfff;
      20'h042da: out <= 12'hfff;
      20'h042db: out <= 12'hfff;
      20'h042dc: out <= 12'hc7f;
      20'h042dd: out <= 12'hc7f;
      20'h042de: out <= 12'h72f;
      20'h042df: out <= 12'h72f;
      20'h042e0: out <= 12'h72f;
      20'h042e1: out <= 12'h72f;
      20'h042e2: out <= 12'h72f;
      20'h042e3: out <= 12'hc7f;
      20'h042e4: out <= 12'hc7f;
      20'h042e5: out <= 12'hfff;
      20'h042e6: out <= 12'hfff;
      20'h042e7: out <= 12'hfff;
      20'h042e8: out <= 12'h222;
      20'h042e9: out <= 12'hfff;
      20'h042ea: out <= 12'hfff;
      20'h042eb: out <= 12'hfff;
      20'h042ec: out <= 12'hc7f;
      20'h042ed: out <= 12'hc7f;
      20'h042ee: out <= 12'hfff;
      20'h042ef: out <= 12'hfff;
      20'h042f0: out <= 12'hfff;
      20'h042f1: out <= 12'hfff;
      20'h042f2: out <= 12'hfff;
      20'h042f3: out <= 12'hc7f;
      20'h042f4: out <= 12'hc7f;
      20'h042f5: out <= 12'hfff;
      20'h042f6: out <= 12'hfff;
      20'h042f7: out <= 12'hfff;
      20'h042f8: out <= 12'h000;
      20'h042f9: out <= 12'h000;
      20'h042fa: out <= 12'h000;
      20'h042fb: out <= 12'h72f;
      20'h042fc: out <= 12'hfff;
      20'h042fd: out <= 12'h72f;
      20'h042fe: out <= 12'hfff;
      20'h042ff: out <= 12'hc7f;
      20'h04300: out <= 12'hc7f;
      20'h04301: out <= 12'hc7f;
      20'h04302: out <= 12'hc7f;
      20'h04303: out <= 12'hc7f;
      20'h04304: out <= 12'hfff;
      20'h04305: out <= 12'hfff;
      20'h04306: out <= 12'h72f;
      20'h04307: out <= 12'h000;
      20'h04308: out <= 12'h222;
      20'h04309: out <= 12'h222;
      20'h0430a: out <= 12'h222;
      20'h0430b: out <= 12'h72f;
      20'h0430c: out <= 12'hfff;
      20'h0430d: out <= 12'h72f;
      20'h0430e: out <= 12'h72f;
      20'h0430f: out <= 12'hc7f;
      20'h04310: out <= 12'hc7f;
      20'h04311: out <= 12'hc7f;
      20'h04312: out <= 12'hc7f;
      20'h04313: out <= 12'hc7f;
      20'h04314: out <= 12'h72f;
      20'h04315: out <= 12'hfff;
      20'h04316: out <= 12'h72f;
      20'h04317: out <= 12'h222;
      20'h04318: out <= 12'h000;
      20'h04319: out <= 12'h000;
      20'h0431a: out <= 12'h000;
      20'h0431b: out <= 12'h000;
      20'h0431c: out <= 12'h000;
      20'h0431d: out <= 12'h000;
      20'h0431e: out <= 12'h000;
      20'h0431f: out <= 12'h72f;
      20'h04320: out <= 12'hfff;
      20'h04321: out <= 12'h72f;
      20'h04322: out <= 12'h000;
      20'h04323: out <= 12'h000;
      20'h04324: out <= 12'h000;
      20'h04325: out <= 12'h000;
      20'h04326: out <= 12'h000;
      20'h04327: out <= 12'h000;
      20'h04328: out <= 12'h222;
      20'h04329: out <= 12'h222;
      20'h0432a: out <= 12'h222;
      20'h0432b: out <= 12'h222;
      20'h0432c: out <= 12'h222;
      20'h0432d: out <= 12'h222;
      20'h0432e: out <= 12'h222;
      20'h0432f: out <= 12'h72f;
      20'h04330: out <= 12'hfff;
      20'h04331: out <= 12'h72f;
      20'h04332: out <= 12'h222;
      20'h04333: out <= 12'h222;
      20'h04334: out <= 12'h222;
      20'h04335: out <= 12'h222;
      20'h04336: out <= 12'h222;
      20'h04337: out <= 12'h222;
      20'h04338: out <= 12'h603;
      20'h04339: out <= 12'h603;
      20'h0433a: out <= 12'h603;
      20'h0433b: out <= 12'h603;
      20'h0433c: out <= 12'h000;
      20'h0433d: out <= 12'h000;
      20'h0433e: out <= 12'hee9;
      20'h0433f: out <= 12'hb27;
      20'h04340: out <= 12'hb27;
      20'h04341: out <= 12'hb27;
      20'h04342: out <= 12'hb27;
      20'h04343: out <= 12'hb27;
      20'h04344: out <= 12'hb27;
      20'h04345: out <= 12'hb27;
      20'h04346: out <= 12'hb27;
      20'h04347: out <= 12'hb27;
      20'h04348: out <= 12'hb27;
      20'h04349: out <= 12'hb27;
      20'h0434a: out <= 12'hee9;
      20'h0434b: out <= 12'h000;
      20'h0434c: out <= 12'h000;
      20'h0434d: out <= 12'hee9;
      20'h0434e: out <= 12'hf87;
      20'h0434f: out <= 12'hf87;
      20'h04350: out <= 12'hb27;
      20'h04351: out <= 12'hee9;
      20'h04352: out <= 12'hee9;
      20'h04353: out <= 12'hee9;
      20'h04354: out <= 12'hee9;
      20'h04355: out <= 12'hee9;
      20'h04356: out <= 12'hee9;
      20'h04357: out <= 12'hee9;
      20'h04358: out <= 12'hb27;
      20'h04359: out <= 12'hf87;
      20'h0435a: out <= 12'hf87;
      20'h0435b: out <= 12'hb27;
      20'h0435c: out <= 12'h000;
      20'h0435d: out <= 12'hee9;
      20'h0435e: out <= 12'hf87;
      20'h0435f: out <= 12'hf87;
      20'h04360: out <= 12'hb27;
      20'h04361: out <= 12'hee9;
      20'h04362: out <= 12'hee9;
      20'h04363: out <= 12'hee9;
      20'h04364: out <= 12'hee9;
      20'h04365: out <= 12'hee9;
      20'h04366: out <= 12'hee9;
      20'h04367: out <= 12'hee9;
      20'h04368: out <= 12'hb27;
      20'h04369: out <= 12'hf87;
      20'h0436a: out <= 12'hf87;
      20'h0436b: out <= 12'hb27;
      20'h0436c: out <= 12'h603;
      20'h0436d: out <= 12'h603;
      20'h0436e: out <= 12'h603;
      20'h0436f: out <= 12'h603;
      20'h04370: out <= 12'h603;
      20'h04371: out <= 12'h603;
      20'h04372: out <= 12'h603;
      20'h04373: out <= 12'h603;
      20'h04374: out <= 12'h603;
      20'h04375: out <= 12'h603;
      20'h04376: out <= 12'h603;
      20'h04377: out <= 12'h603;
      20'h04378: out <= 12'h603;
      20'h04379: out <= 12'h603;
      20'h0437a: out <= 12'h603;
      20'h0437b: out <= 12'h603;
      20'h0437c: out <= 12'h603;
      20'h0437d: out <= 12'h603;
      20'h0437e: out <= 12'h603;
      20'h0437f: out <= 12'h603;
      20'h04380: out <= 12'h603;
      20'h04381: out <= 12'h603;
      20'h04382: out <= 12'h603;
      20'h04383: out <= 12'h603;
      20'h04384: out <= 12'h603;
      20'h04385: out <= 12'h603;
      20'h04386: out <= 12'h603;
      20'h04387: out <= 12'h603;
      20'h04388: out <= 12'h603;
      20'h04389: out <= 12'h603;
      20'h0438a: out <= 12'h603;
      20'h0438b: out <= 12'h603;
      20'h0438c: out <= 12'h603;
      20'h0438d: out <= 12'h603;
      20'h0438e: out <= 12'h603;
      20'h0438f: out <= 12'h603;
      20'h04390: out <= 12'hee9;
      20'h04391: out <= 12'hf87;
      20'h04392: out <= 12'hee9;
      20'h04393: out <= 12'hb27;
      20'h04394: out <= 12'hb27;
      20'h04395: out <= 12'hb27;
      20'h04396: out <= 12'hf87;
      20'h04397: out <= 12'hb27;
      20'h04398: out <= 12'h000;
      20'h04399: out <= 12'h000;
      20'h0439a: out <= 12'h000;
      20'h0439b: out <= 12'h000;
      20'h0439c: out <= 12'h000;
      20'h0439d: out <= 12'h000;
      20'h0439e: out <= 12'h000;
      20'h0439f: out <= 12'h000;
      20'h043a0: out <= 12'h000;
      20'h043a1: out <= 12'h000;
      20'h043a2: out <= 12'h000;
      20'h043a3: out <= 12'h000;
      20'h043a4: out <= 12'h000;
      20'h043a5: out <= 12'h000;
      20'h043a6: out <= 12'h000;
      20'h043a7: out <= 12'h000;
      20'h043a8: out <= 12'h000;
      20'h043a9: out <= 12'h000;
      20'h043aa: out <= 12'h000;
      20'h043ab: out <= 12'h000;
      20'h043ac: out <= 12'h000;
      20'h043ad: out <= 12'h000;
      20'h043ae: out <= 12'h000;
      20'h043af: out <= 12'h000;
      20'h043b0: out <= 12'h000;
      20'h043b1: out <= 12'h000;
      20'h043b2: out <= 12'h000;
      20'h043b3: out <= 12'h000;
      20'h043b4: out <= 12'h000;
      20'h043b5: out <= 12'h000;
      20'h043b6: out <= 12'h000;
      20'h043b7: out <= 12'h000;
      20'h043b8: out <= 12'h000;
      20'h043b9: out <= 12'h000;
      20'h043ba: out <= 12'h000;
      20'h043bb: out <= 12'h000;
      20'h043bc: out <= 12'h000;
      20'h043bd: out <= 12'h000;
      20'h043be: out <= 12'h000;
      20'h043bf: out <= 12'h000;
      20'h043c0: out <= 12'h000;
      20'h043c1: out <= 12'h000;
      20'h043c2: out <= 12'h000;
      20'h043c3: out <= 12'h000;
      20'h043c4: out <= 12'h000;
      20'h043c5: out <= 12'h000;
      20'h043c6: out <= 12'h000;
      20'h043c7: out <= 12'h000;
      20'h043c8: out <= 12'h000;
      20'h043c9: out <= 12'h000;
      20'h043ca: out <= 12'h000;
      20'h043cb: out <= 12'h000;
      20'h043cc: out <= 12'h000;
      20'h043cd: out <= 12'h000;
      20'h043ce: out <= 12'h000;
      20'h043cf: out <= 12'h000;
      20'h043d0: out <= 12'h000;
      20'h043d1: out <= 12'hc7f;
      20'h043d2: out <= 12'hfff;
      20'h043d3: out <= 12'hc7f;
      20'h043d4: out <= 12'hfff;
      20'h043d5: out <= 12'hfff;
      20'h043d6: out <= 12'hfff;
      20'h043d7: out <= 12'hfff;
      20'h043d8: out <= 12'hfff;
      20'h043d9: out <= 12'hc7f;
      20'h043da: out <= 12'hc7f;
      20'h043db: out <= 12'hfff;
      20'h043dc: out <= 12'hc7f;
      20'h043dd: out <= 12'h000;
      20'h043de: out <= 12'h000;
      20'h043df: out <= 12'h000;
      20'h043e0: out <= 12'h222;
      20'h043e1: out <= 12'hc7f;
      20'h043e2: out <= 12'hfff;
      20'h043e3: out <= 12'hc7f;
      20'h043e4: out <= 12'h72f;
      20'h043e5: out <= 12'h72f;
      20'h043e6: out <= 12'h72f;
      20'h043e7: out <= 12'h72f;
      20'h043e8: out <= 12'h72f;
      20'h043e9: out <= 12'hc7f;
      20'h043ea: out <= 12'hc7f;
      20'h043eb: out <= 12'hfff;
      20'h043ec: out <= 12'hc7f;
      20'h043ed: out <= 12'h222;
      20'h043ee: out <= 12'h222;
      20'h043ef: out <= 12'h222;
      20'h043f0: out <= 12'h000;
      20'h043f1: out <= 12'hc7f;
      20'h043f2: out <= 12'h72f;
      20'h043f3: out <= 12'hc7f;
      20'h043f4: out <= 12'hfff;
      20'h043f5: out <= 12'hfff;
      20'h043f6: out <= 12'hc7f;
      20'h043f7: out <= 12'hc7f;
      20'h043f8: out <= 12'hc7f;
      20'h043f9: out <= 12'hc7f;
      20'h043fa: out <= 12'hc7f;
      20'h043fb: out <= 12'hfff;
      20'h043fc: out <= 12'hfff;
      20'h043fd: out <= 12'hc7f;
      20'h043fe: out <= 12'h72f;
      20'h043ff: out <= 12'hc7f;
      20'h04400: out <= 12'h222;
      20'h04401: out <= 12'hc7f;
      20'h04402: out <= 12'h72f;
      20'h04403: out <= 12'hc7f;
      20'h04404: out <= 12'h72f;
      20'h04405: out <= 12'h72f;
      20'h04406: out <= 12'hc7f;
      20'h04407: out <= 12'hc7f;
      20'h04408: out <= 12'hc7f;
      20'h04409: out <= 12'hc7f;
      20'h0440a: out <= 12'hc7f;
      20'h0440b: out <= 12'h72f;
      20'h0440c: out <= 12'h72f;
      20'h0440d: out <= 12'hc7f;
      20'h0440e: out <= 12'h72f;
      20'h0440f: out <= 12'hc7f;
      20'h04410: out <= 12'h000;
      20'h04411: out <= 12'h000;
      20'h04412: out <= 12'h000;
      20'h04413: out <= 12'hc7f;
      20'h04414: out <= 12'hfff;
      20'h04415: out <= 12'hc7f;
      20'h04416: out <= 12'hc7f;
      20'h04417: out <= 12'hfff;
      20'h04418: out <= 12'hfff;
      20'h04419: out <= 12'hfff;
      20'h0441a: out <= 12'hfff;
      20'h0441b: out <= 12'hfff;
      20'h0441c: out <= 12'hc7f;
      20'h0441d: out <= 12'hfff;
      20'h0441e: out <= 12'hc7f;
      20'h0441f: out <= 12'h000;
      20'h04420: out <= 12'h222;
      20'h04421: out <= 12'h222;
      20'h04422: out <= 12'h222;
      20'h04423: out <= 12'hc7f;
      20'h04424: out <= 12'hfff;
      20'h04425: out <= 12'hc7f;
      20'h04426: out <= 12'hc7f;
      20'h04427: out <= 12'h72f;
      20'h04428: out <= 12'h72f;
      20'h04429: out <= 12'h72f;
      20'h0442a: out <= 12'h72f;
      20'h0442b: out <= 12'h72f;
      20'h0442c: out <= 12'hc7f;
      20'h0442d: out <= 12'hfff;
      20'h0442e: out <= 12'hc7f;
      20'h0442f: out <= 12'h222;
      20'h04430: out <= 12'h000;
      20'h04431: out <= 12'h000;
      20'h04432: out <= 12'h000;
      20'h04433: out <= 12'h000;
      20'h04434: out <= 12'h000;
      20'h04435: out <= 12'h000;
      20'h04436: out <= 12'h000;
      20'h04437: out <= 12'h72f;
      20'h04438: out <= 12'hfff;
      20'h04439: out <= 12'h72f;
      20'h0443a: out <= 12'h000;
      20'h0443b: out <= 12'h000;
      20'h0443c: out <= 12'h000;
      20'h0443d: out <= 12'h000;
      20'h0443e: out <= 12'h000;
      20'h0443f: out <= 12'h000;
      20'h04440: out <= 12'h222;
      20'h04441: out <= 12'h222;
      20'h04442: out <= 12'h222;
      20'h04443: out <= 12'h222;
      20'h04444: out <= 12'h222;
      20'h04445: out <= 12'h222;
      20'h04446: out <= 12'h222;
      20'h04447: out <= 12'h72f;
      20'h04448: out <= 12'hfff;
      20'h04449: out <= 12'h72f;
      20'h0444a: out <= 12'h222;
      20'h0444b: out <= 12'h222;
      20'h0444c: out <= 12'h222;
      20'h0444d: out <= 12'h222;
      20'h0444e: out <= 12'h222;
      20'h0444f: out <= 12'h222;
      20'h04450: out <= 12'h603;
      20'h04451: out <= 12'h603;
      20'h04452: out <= 12'h603;
      20'h04453: out <= 12'h603;
      20'h04454: out <= 12'h000;
      20'h04455: out <= 12'h000;
      20'h04456: out <= 12'h000;
      20'h04457: out <= 12'h000;
      20'h04458: out <= 12'h000;
      20'h04459: out <= 12'h000;
      20'h0445a: out <= 12'h000;
      20'h0445b: out <= 12'h000;
      20'h0445c: out <= 12'h000;
      20'h0445d: out <= 12'h000;
      20'h0445e: out <= 12'h000;
      20'h0445f: out <= 12'h000;
      20'h04460: out <= 12'h000;
      20'h04461: out <= 12'h000;
      20'h04462: out <= 12'h000;
      20'h04463: out <= 12'h000;
      20'h04464: out <= 12'h000;
      20'h04465: out <= 12'hee9;
      20'h04466: out <= 12'hb27;
      20'h04467: out <= 12'hb27;
      20'h04468: out <= 12'hf87;
      20'h04469: out <= 12'hf87;
      20'h0446a: out <= 12'hf87;
      20'h0446b: out <= 12'hf87;
      20'h0446c: out <= 12'hf87;
      20'h0446d: out <= 12'hf87;
      20'h0446e: out <= 12'hf87;
      20'h0446f: out <= 12'hf87;
      20'h04470: out <= 12'hf87;
      20'h04471: out <= 12'hb27;
      20'h04472: out <= 12'hb27;
      20'h04473: out <= 12'hb27;
      20'h04474: out <= 12'h000;
      20'h04475: out <= 12'hee9;
      20'h04476: out <= 12'hb27;
      20'h04477: out <= 12'hb27;
      20'h04478: out <= 12'hf87;
      20'h04479: out <= 12'hf87;
      20'h0447a: out <= 12'hf87;
      20'h0447b: out <= 12'hf87;
      20'h0447c: out <= 12'hf87;
      20'h0447d: out <= 12'hf87;
      20'h0447e: out <= 12'hf87;
      20'h0447f: out <= 12'hf87;
      20'h04480: out <= 12'hf87;
      20'h04481: out <= 12'hb27;
      20'h04482: out <= 12'hb27;
      20'h04483: out <= 12'hb27;
      20'h04484: out <= 12'h603;
      20'h04485: out <= 12'h603;
      20'h04486: out <= 12'h603;
      20'h04487: out <= 12'h603;
      20'h04488: out <= 12'h603;
      20'h04489: out <= 12'h603;
      20'h0448a: out <= 12'h603;
      20'h0448b: out <= 12'h603;
      20'h0448c: out <= 12'h603;
      20'h0448d: out <= 12'h603;
      20'h0448e: out <= 12'h603;
      20'h0448f: out <= 12'h603;
      20'h04490: out <= 12'h603;
      20'h04491: out <= 12'h603;
      20'h04492: out <= 12'h603;
      20'h04493: out <= 12'h603;
      20'h04494: out <= 12'h603;
      20'h04495: out <= 12'h603;
      20'h04496: out <= 12'h603;
      20'h04497: out <= 12'h603;
      20'h04498: out <= 12'h603;
      20'h04499: out <= 12'h603;
      20'h0449a: out <= 12'h603;
      20'h0449b: out <= 12'h603;
      20'h0449c: out <= 12'h603;
      20'h0449d: out <= 12'h603;
      20'h0449e: out <= 12'h603;
      20'h0449f: out <= 12'h603;
      20'h044a0: out <= 12'h603;
      20'h044a1: out <= 12'h603;
      20'h044a2: out <= 12'h603;
      20'h044a3: out <= 12'h603;
      20'h044a4: out <= 12'h603;
      20'h044a5: out <= 12'h603;
      20'h044a6: out <= 12'h603;
      20'h044a7: out <= 12'h603;
      20'h044a8: out <= 12'hee9;
      20'h044a9: out <= 12'hf87;
      20'h044aa: out <= 12'hf87;
      20'h044ab: out <= 12'hf87;
      20'h044ac: out <= 12'hf87;
      20'h044ad: out <= 12'hf87;
      20'h044ae: out <= 12'hf87;
      20'h044af: out <= 12'hb27;
      20'h044b0: out <= 12'h000;
      20'h044b1: out <= 12'h000;
      20'h044b2: out <= 12'h000;
      20'h044b3: out <= 12'h000;
      20'h044b4: out <= 12'h000;
      20'h044b5: out <= 12'h000;
      20'h044b6: out <= 12'h000;
      20'h044b7: out <= 12'h000;
      20'h044b8: out <= 12'h000;
      20'h044b9: out <= 12'h000;
      20'h044ba: out <= 12'h000;
      20'h044bb: out <= 12'h000;
      20'h044bc: out <= 12'h000;
      20'h044bd: out <= 12'h000;
      20'h044be: out <= 12'h000;
      20'h044bf: out <= 12'h000;
      20'h044c0: out <= 12'h000;
      20'h044c1: out <= 12'h000;
      20'h044c2: out <= 12'h000;
      20'h044c3: out <= 12'h000;
      20'h044c4: out <= 12'h000;
      20'h044c5: out <= 12'h000;
      20'h044c6: out <= 12'h000;
      20'h044c7: out <= 12'h000;
      20'h044c8: out <= 12'h000;
      20'h044c9: out <= 12'h000;
      20'h044ca: out <= 12'h000;
      20'h044cb: out <= 12'h000;
      20'h044cc: out <= 12'h000;
      20'h044cd: out <= 12'h000;
      20'h044ce: out <= 12'h000;
      20'h044cf: out <= 12'h000;
      20'h044d0: out <= 12'h000;
      20'h044d1: out <= 12'h000;
      20'h044d2: out <= 12'h000;
      20'h044d3: out <= 12'h000;
      20'h044d4: out <= 12'h000;
      20'h044d5: out <= 12'h000;
      20'h044d6: out <= 12'h000;
      20'h044d7: out <= 12'h000;
      20'h044d8: out <= 12'h000;
      20'h044d9: out <= 12'h000;
      20'h044da: out <= 12'h000;
      20'h044db: out <= 12'h000;
      20'h044dc: out <= 12'h000;
      20'h044dd: out <= 12'h000;
      20'h044de: out <= 12'h000;
      20'h044df: out <= 12'h000;
      20'h044e0: out <= 12'h000;
      20'h044e1: out <= 12'h000;
      20'h044e2: out <= 12'h000;
      20'h044e3: out <= 12'h000;
      20'h044e4: out <= 12'h000;
      20'h044e5: out <= 12'h000;
      20'h044e6: out <= 12'h000;
      20'h044e7: out <= 12'h000;
      20'h044e8: out <= 12'h000;
      20'h044e9: out <= 12'h000;
      20'h044ea: out <= 12'h000;
      20'h044eb: out <= 12'h000;
      20'h044ec: out <= 12'h000;
      20'h044ed: out <= 12'h000;
      20'h044ee: out <= 12'h000;
      20'h044ef: out <= 12'h000;
      20'h044f0: out <= 12'h000;
      20'h044f1: out <= 12'h000;
      20'h044f2: out <= 12'h000;
      20'h044f3: out <= 12'h000;
      20'h044f4: out <= 12'h000;
      20'h044f5: out <= 12'h000;
      20'h044f6: out <= 12'h000;
      20'h044f7: out <= 12'h000;
      20'h044f8: out <= 12'h222;
      20'h044f9: out <= 12'h222;
      20'h044fa: out <= 12'h222;
      20'h044fb: out <= 12'h222;
      20'h044fc: out <= 12'h222;
      20'h044fd: out <= 12'h222;
      20'h044fe: out <= 12'h222;
      20'h044ff: out <= 12'h222;
      20'h04500: out <= 12'h222;
      20'h04501: out <= 12'h222;
      20'h04502: out <= 12'h222;
      20'h04503: out <= 12'h222;
      20'h04504: out <= 12'h222;
      20'h04505: out <= 12'h222;
      20'h04506: out <= 12'h222;
      20'h04507: out <= 12'h222;
      20'h04508: out <= 12'h000;
      20'h04509: out <= 12'h000;
      20'h0450a: out <= 12'h000;
      20'h0450b: out <= 12'h000;
      20'h0450c: out <= 12'h000;
      20'h0450d: out <= 12'h000;
      20'h0450e: out <= 12'hfff;
      20'h0450f: out <= 12'hfff;
      20'h04510: out <= 12'hfff;
      20'h04511: out <= 12'hfff;
      20'h04512: out <= 12'hfff;
      20'h04513: out <= 12'h000;
      20'h04514: out <= 12'h000;
      20'h04515: out <= 12'h000;
      20'h04516: out <= 12'h000;
      20'h04517: out <= 12'h000;
      20'h04518: out <= 12'h222;
      20'h04519: out <= 12'h222;
      20'h0451a: out <= 12'h222;
      20'h0451b: out <= 12'h222;
      20'h0451c: out <= 12'h222;
      20'h0451d: out <= 12'h222;
      20'h0451e: out <= 12'h72f;
      20'h0451f: out <= 12'h72f;
      20'h04520: out <= 12'h72f;
      20'h04521: out <= 12'h72f;
      20'h04522: out <= 12'h72f;
      20'h04523: out <= 12'h222;
      20'h04524: out <= 12'h222;
      20'h04525: out <= 12'h222;
      20'h04526: out <= 12'h222;
      20'h04527: out <= 12'h222;
      20'h04528: out <= 12'h000;
      20'h04529: out <= 12'h000;
      20'h0452a: out <= 12'h000;
      20'h0452b: out <= 12'h000;
      20'h0452c: out <= 12'h000;
      20'h0452d: out <= 12'h000;
      20'h0452e: out <= 12'h000;
      20'h0452f: out <= 12'h000;
      20'h04530: out <= 12'h000;
      20'h04531: out <= 12'h000;
      20'h04532: out <= 12'h000;
      20'h04533: out <= 12'h000;
      20'h04534: out <= 12'h000;
      20'h04535: out <= 12'h000;
      20'h04536: out <= 12'h000;
      20'h04537: out <= 12'h000;
      20'h04538: out <= 12'h222;
      20'h04539: out <= 12'h222;
      20'h0453a: out <= 12'h222;
      20'h0453b: out <= 12'h222;
      20'h0453c: out <= 12'h222;
      20'h0453d: out <= 12'h222;
      20'h0453e: out <= 12'h222;
      20'h0453f: out <= 12'h222;
      20'h04540: out <= 12'h222;
      20'h04541: out <= 12'h222;
      20'h04542: out <= 12'h222;
      20'h04543: out <= 12'h222;
      20'h04544: out <= 12'h222;
      20'h04545: out <= 12'h222;
      20'h04546: out <= 12'h222;
      20'h04547: out <= 12'h222;
      20'h04548: out <= 12'h000;
      20'h04549: out <= 12'h000;
      20'h0454a: out <= 12'h000;
      20'h0454b: out <= 12'h000;
      20'h0454c: out <= 12'h000;
      20'h0454d: out <= 12'h000;
      20'h0454e: out <= 12'h000;
      20'h0454f: out <= 12'hc7f;
      20'h04550: out <= 12'hfff;
      20'h04551: out <= 12'hc7f;
      20'h04552: out <= 12'h000;
      20'h04553: out <= 12'h000;
      20'h04554: out <= 12'h000;
      20'h04555: out <= 12'h000;
      20'h04556: out <= 12'h000;
      20'h04557: out <= 12'h000;
      20'h04558: out <= 12'h222;
      20'h04559: out <= 12'h222;
      20'h0455a: out <= 12'h222;
      20'h0455b: out <= 12'h222;
      20'h0455c: out <= 12'h222;
      20'h0455d: out <= 12'h222;
      20'h0455e: out <= 12'h222;
      20'h0455f: out <= 12'hc7f;
      20'h04560: out <= 12'hfff;
      20'h04561: out <= 12'hc7f;
      20'h04562: out <= 12'h222;
      20'h04563: out <= 12'h222;
      20'h04564: out <= 12'h222;
      20'h04565: out <= 12'h222;
      20'h04566: out <= 12'h222;
      20'h04567: out <= 12'h222;
      20'h04568: out <= 12'h603;
      20'h04569: out <= 12'h603;
      20'h0456a: out <= 12'h603;
      20'h0456b: out <= 12'h603;
      20'h0456c: out <= 12'h000;
      20'h0456d: out <= 12'h000;
      20'h0456e: out <= 12'h000;
      20'h0456f: out <= 12'h000;
      20'h04570: out <= 12'h000;
      20'h04571: out <= 12'h000;
      20'h04572: out <= 12'h000;
      20'h04573: out <= 12'h000;
      20'h04574: out <= 12'h000;
      20'h04575: out <= 12'h000;
      20'h04576: out <= 12'h000;
      20'h04577: out <= 12'h000;
      20'h04578: out <= 12'h000;
      20'h04579: out <= 12'h000;
      20'h0457a: out <= 12'h000;
      20'h0457b: out <= 12'h000;
      20'h0457c: out <= 12'h000;
      20'h0457d: out <= 12'h000;
      20'h0457e: out <= 12'h000;
      20'h0457f: out <= 12'h000;
      20'h04580: out <= 12'h000;
      20'h04581: out <= 12'h000;
      20'h04582: out <= 12'h000;
      20'h04583: out <= 12'h000;
      20'h04584: out <= 12'h000;
      20'h04585: out <= 12'h000;
      20'h04586: out <= 12'h000;
      20'h04587: out <= 12'h000;
      20'h04588: out <= 12'h000;
      20'h04589: out <= 12'h000;
      20'h0458a: out <= 12'h000;
      20'h0458b: out <= 12'h000;
      20'h0458c: out <= 12'h000;
      20'h0458d: out <= 12'h000;
      20'h0458e: out <= 12'h000;
      20'h0458f: out <= 12'h000;
      20'h04590: out <= 12'h000;
      20'h04591: out <= 12'h000;
      20'h04592: out <= 12'h000;
      20'h04593: out <= 12'h000;
      20'h04594: out <= 12'h000;
      20'h04595: out <= 12'h000;
      20'h04596: out <= 12'h000;
      20'h04597: out <= 12'h000;
      20'h04598: out <= 12'h000;
      20'h04599: out <= 12'h000;
      20'h0459a: out <= 12'h000;
      20'h0459b: out <= 12'h000;
      20'h0459c: out <= 12'h603;
      20'h0459d: out <= 12'h603;
      20'h0459e: out <= 12'h603;
      20'h0459f: out <= 12'h603;
      20'h045a0: out <= 12'h603;
      20'h045a1: out <= 12'h603;
      20'h045a2: out <= 12'h603;
      20'h045a3: out <= 12'h603;
      20'h045a4: out <= 12'h603;
      20'h045a5: out <= 12'h603;
      20'h045a6: out <= 12'h603;
      20'h045a7: out <= 12'h603;
      20'h045a8: out <= 12'h603;
      20'h045a9: out <= 12'h603;
      20'h045aa: out <= 12'h603;
      20'h045ab: out <= 12'h603;
      20'h045ac: out <= 12'h603;
      20'h045ad: out <= 12'h603;
      20'h045ae: out <= 12'h603;
      20'h045af: out <= 12'h603;
      20'h045b0: out <= 12'h603;
      20'h045b1: out <= 12'h603;
      20'h045b2: out <= 12'h603;
      20'h045b3: out <= 12'h603;
      20'h045b4: out <= 12'h603;
      20'h045b5: out <= 12'h603;
      20'h045b6: out <= 12'h603;
      20'h045b7: out <= 12'h603;
      20'h045b8: out <= 12'h603;
      20'h045b9: out <= 12'h603;
      20'h045ba: out <= 12'h603;
      20'h045bb: out <= 12'h603;
      20'h045bc: out <= 12'h603;
      20'h045bd: out <= 12'h603;
      20'h045be: out <= 12'h603;
      20'h045bf: out <= 12'h603;
      20'h045c0: out <= 12'hb27;
      20'h045c1: out <= 12'hb27;
      20'h045c2: out <= 12'hb27;
      20'h045c3: out <= 12'hb27;
      20'h045c4: out <= 12'hb27;
      20'h045c5: out <= 12'hb27;
      20'h045c6: out <= 12'hb27;
      20'h045c7: out <= 12'hb27;
      20'h045c8: out <= 12'h000;
      20'h045c9: out <= 12'h000;
      20'h045ca: out <= 12'h000;
      20'h045cb: out <= 12'h000;
      20'h045cc: out <= 12'h000;
      20'h045cd: out <= 12'h000;
      20'h045ce: out <= 12'h000;
      20'h045cf: out <= 12'h000;
      20'h045d0: out <= 12'h000;
      20'h045d1: out <= 12'h000;
      20'h045d2: out <= 12'h000;
      20'h045d3: out <= 12'h000;
      20'h045d4: out <= 12'h000;
      20'h045d5: out <= 12'h000;
      20'h045d6: out <= 12'h000;
      20'h045d7: out <= 12'h000;
      20'h045d8: out <= 12'h000;
      20'h045d9: out <= 12'h000;
      20'h045da: out <= 12'h000;
      20'h045db: out <= 12'h000;
      20'h045dc: out <= 12'h000;
      20'h045dd: out <= 12'h000;
      20'h045de: out <= 12'h000;
      20'h045df: out <= 12'h000;
      20'h045e0: out <= 12'h000;
      20'h045e1: out <= 12'h000;
      20'h045e2: out <= 12'h000;
      20'h045e3: out <= 12'h000;
      20'h045e4: out <= 12'h000;
      20'h045e5: out <= 12'h000;
      20'h045e6: out <= 12'h000;
      20'h045e7: out <= 12'h000;
      20'h045e8: out <= 12'h000;
      20'h045e9: out <= 12'h000;
      20'h045ea: out <= 12'h000;
      20'h045eb: out <= 12'h000;
      20'h045ec: out <= 12'h000;
      20'h045ed: out <= 12'h000;
      20'h045ee: out <= 12'h000;
      20'h045ef: out <= 12'h000;
      20'h045f0: out <= 12'h000;
      20'h045f1: out <= 12'h000;
      20'h045f2: out <= 12'h000;
      20'h045f3: out <= 12'h000;
      20'h045f4: out <= 12'h000;
      20'h045f5: out <= 12'h000;
      20'h045f6: out <= 12'h000;
      20'h045f7: out <= 12'h000;
      20'h045f8: out <= 12'h000;
      20'h045f9: out <= 12'h000;
      20'h045fa: out <= 12'h000;
      20'h045fb: out <= 12'h000;
      20'h045fc: out <= 12'h000;
      20'h045fd: out <= 12'h000;
      20'h045fe: out <= 12'h000;
      20'h045ff: out <= 12'h000;
      20'h04600: out <= 12'h603;
      20'h04601: out <= 12'h603;
      20'h04602: out <= 12'h603;
      20'h04603: out <= 12'h603;
      20'h04604: out <= 12'h603;
      20'h04605: out <= 12'h603;
      20'h04606: out <= 12'h603;
      20'h04607: out <= 12'h603;
      20'h04608: out <= 12'h603;
      20'h04609: out <= 12'h603;
      20'h0460a: out <= 12'h603;
      20'h0460b: out <= 12'h603;
      20'h0460c: out <= 12'h603;
      20'h0460d: out <= 12'h603;
      20'h0460e: out <= 12'h603;
      20'h0460f: out <= 12'h603;
      20'h04610: out <= 12'h603;
      20'h04611: out <= 12'h603;
      20'h04612: out <= 12'h603;
      20'h04613: out <= 12'h603;
      20'h04614: out <= 12'h603;
      20'h04615: out <= 12'h603;
      20'h04616: out <= 12'h603;
      20'h04617: out <= 12'h603;
      20'h04618: out <= 12'h603;
      20'h04619: out <= 12'h603;
      20'h0461a: out <= 12'h603;
      20'h0461b: out <= 12'h603;
      20'h0461c: out <= 12'h603;
      20'h0461d: out <= 12'h603;
      20'h0461e: out <= 12'h603;
      20'h0461f: out <= 12'h603;
      20'h04620: out <= 12'h603;
      20'h04621: out <= 12'h603;
      20'h04622: out <= 12'h603;
      20'h04623: out <= 12'h603;
      20'h04624: out <= 12'h603;
      20'h04625: out <= 12'h603;
      20'h04626: out <= 12'h603;
      20'h04627: out <= 12'h603;
      20'h04628: out <= 12'h603;
      20'h04629: out <= 12'h603;
      20'h0462a: out <= 12'h603;
      20'h0462b: out <= 12'h603;
      20'h0462c: out <= 12'h603;
      20'h0462d: out <= 12'h603;
      20'h0462e: out <= 12'h603;
      20'h0462f: out <= 12'h603;
      20'h04630: out <= 12'h603;
      20'h04631: out <= 12'h603;
      20'h04632: out <= 12'h603;
      20'h04633: out <= 12'h603;
      20'h04634: out <= 12'h000;
      20'h04635: out <= 12'h000;
      20'h04636: out <= 12'h000;
      20'h04637: out <= 12'h6af;
      20'h04638: out <= 12'hfff;
      20'h04639: out <= 12'h6af;
      20'h0463a: out <= 12'h000;
      20'h0463b: out <= 12'h000;
      20'h0463c: out <= 12'h603;
      20'h0463d: out <= 12'h603;
      20'h0463e: out <= 12'h603;
      20'h0463f: out <= 12'h603;
      20'h04640: out <= 12'h603;
      20'h04641: out <= 12'h603;
      20'h04642: out <= 12'h603;
      20'h04643: out <= 12'h603;
      20'h04644: out <= 12'h603;
      20'h04645: out <= 12'h603;
      20'h04646: out <= 12'h603;
      20'h04647: out <= 12'h603;
      20'h04648: out <= 12'h603;
      20'h04649: out <= 12'h603;
      20'h0464a: out <= 12'h603;
      20'h0464b: out <= 12'h603;
      20'h0464c: out <= 12'h603;
      20'h0464d: out <= 12'h603;
      20'h0464e: out <= 12'h603;
      20'h0464f: out <= 12'h603;
      20'h04650: out <= 12'h603;
      20'h04651: out <= 12'h603;
      20'h04652: out <= 12'h603;
      20'h04653: out <= 12'h603;
      20'h04654: out <= 12'h000;
      20'h04655: out <= 12'h000;
      20'h04656: out <= 12'h000;
      20'h04657: out <= 12'h660;
      20'h04658: out <= 12'hbb0;
      20'h04659: out <= 12'h660;
      20'h0465a: out <= 12'h000;
      20'h0465b: out <= 12'h000;
      20'h0465c: out <= 12'h603;
      20'h0465d: out <= 12'h603;
      20'h0465e: out <= 12'h603;
      20'h0465f: out <= 12'h603;
      20'h04660: out <= 12'h222;
      20'h04661: out <= 12'h222;
      20'h04662: out <= 12'h222;
      20'h04663: out <= 12'h222;
      20'h04664: out <= 12'h222;
      20'h04665: out <= 12'h222;
      20'h04666: out <= 12'h222;
      20'h04667: out <= 12'h222;
      20'h04668: out <= 12'h222;
      20'h04669: out <= 12'h222;
      20'h0466a: out <= 12'h222;
      20'h0466b: out <= 12'h222;
      20'h0466c: out <= 12'h222;
      20'h0466d: out <= 12'h222;
      20'h0466e: out <= 12'h222;
      20'h0466f: out <= 12'h222;
      20'h04670: out <= 12'h000;
      20'h04671: out <= 12'h000;
      20'h04672: out <= 12'h000;
      20'h04673: out <= 12'h000;
      20'h04674: out <= 12'h000;
      20'h04675: out <= 12'h000;
      20'h04676: out <= 12'h000;
      20'h04677: out <= 12'h000;
      20'h04678: out <= 12'h660;
      20'h04679: out <= 12'h000;
      20'h0467a: out <= 12'h000;
      20'h0467b: out <= 12'h000;
      20'h0467c: out <= 12'h000;
      20'h0467d: out <= 12'h000;
      20'h0467e: out <= 12'h000;
      20'h0467f: out <= 12'h000;
      20'h04680: out <= 12'h603;
      20'h04681: out <= 12'h603;
      20'h04682: out <= 12'h603;
      20'h04683: out <= 12'h603;
      20'h04684: out <= 12'h000;
      20'h04685: out <= 12'h666;
      20'h04686: out <= 12'h666;
      20'h04687: out <= 12'h666;
      20'h04688: out <= 12'h666;
      20'h04689: out <= 12'h666;
      20'h0468a: out <= 12'h666;
      20'h0468b: out <= 12'h666;
      20'h0468c: out <= 12'h666;
      20'h0468d: out <= 12'h666;
      20'h0468e: out <= 12'h666;
      20'h0468f: out <= 12'h666;
      20'h04690: out <= 12'h666;
      20'h04691: out <= 12'h666;
      20'h04692: out <= 12'h666;
      20'h04693: out <= 12'h666;
      20'h04694: out <= 12'h000;
      20'h04695: out <= 12'h000;
      20'h04696: out <= 12'hb27;
      20'h04697: out <= 12'hf87;
      20'h04698: out <= 12'hee9;
      20'h04699: out <= 12'hee9;
      20'h0469a: out <= 12'hf87;
      20'h0469b: out <= 12'hf87;
      20'h0469c: out <= 12'hf87;
      20'h0469d: out <= 12'hf87;
      20'h0469e: out <= 12'hf87;
      20'h0469f: out <= 12'hb27;
      20'h046a0: out <= 12'hb27;
      20'h046a1: out <= 12'hf87;
      20'h046a2: out <= 12'hee9;
      20'h046a3: out <= 12'h000;
      20'h046a4: out <= 12'h000;
      20'h046a5: out <= 12'h000;
      20'h046a6: out <= 12'h000;
      20'h046a7: out <= 12'h000;
      20'h046a8: out <= 12'h000;
      20'h046a9: out <= 12'h000;
      20'h046aa: out <= 12'h000;
      20'h046ab: out <= 12'hee9;
      20'h046ac: out <= 12'hee9;
      20'h046ad: out <= 12'h000;
      20'h046ae: out <= 12'h000;
      20'h046af: out <= 12'h000;
      20'h046b0: out <= 12'h000;
      20'h046b1: out <= 12'h000;
      20'h046b2: out <= 12'h000;
      20'h046b3: out <= 12'h000;
      20'h046b4: out <= 12'h603;
      20'h046b5: out <= 12'h603;
      20'h046b6: out <= 12'h603;
      20'h046b7: out <= 12'h603;
      20'h046b8: out <= 12'h603;
      20'h046b9: out <= 12'h603;
      20'h046ba: out <= 12'h603;
      20'h046bb: out <= 12'h603;
      20'h046bc: out <= 12'h603;
      20'h046bd: out <= 12'h603;
      20'h046be: out <= 12'h603;
      20'h046bf: out <= 12'h603;
      20'h046c0: out <= 12'h603;
      20'h046c1: out <= 12'h603;
      20'h046c2: out <= 12'h603;
      20'h046c3: out <= 12'h603;
      20'h046c4: out <= 12'h603;
      20'h046c5: out <= 12'h603;
      20'h046c6: out <= 12'h603;
      20'h046c7: out <= 12'h603;
      20'h046c8: out <= 12'h603;
      20'h046c9: out <= 12'h603;
      20'h046ca: out <= 12'h603;
      20'h046cb: out <= 12'h603;
      20'h046cc: out <= 12'h603;
      20'h046cd: out <= 12'h603;
      20'h046ce: out <= 12'h603;
      20'h046cf: out <= 12'h603;
      20'h046d0: out <= 12'h603;
      20'h046d1: out <= 12'h603;
      20'h046d2: out <= 12'h603;
      20'h046d3: out <= 12'h603;
      20'h046d4: out <= 12'h603;
      20'h046d5: out <= 12'h603;
      20'h046d6: out <= 12'h603;
      20'h046d7: out <= 12'h603;
      20'h046d8: out <= 12'hee9;
      20'h046d9: out <= 12'hee9;
      20'h046da: out <= 12'hee9;
      20'h046db: out <= 12'hee9;
      20'h046dc: out <= 12'hee9;
      20'h046dd: out <= 12'hee9;
      20'h046de: out <= 12'hee9;
      20'h046df: out <= 12'hb27;
      20'h046e0: out <= 12'h000;
      20'h046e1: out <= 12'h000;
      20'h046e2: out <= 12'h000;
      20'h046e3: out <= 12'h000;
      20'h046e4: out <= 12'h000;
      20'h046e5: out <= 12'h000;
      20'h046e6: out <= 12'h000;
      20'h046e7: out <= 12'h000;
      20'h046e8: out <= 12'h000;
      20'h046e9: out <= 12'h000;
      20'h046ea: out <= 12'h000;
      20'h046eb: out <= 12'h8d0;
      20'h046ec: out <= 12'h8d0;
      20'h046ed: out <= 12'h000;
      20'h046ee: out <= 12'h000;
      20'h046ef: out <= 12'h000;
      20'h046f0: out <= 12'h8d0;
      20'h046f1: out <= 12'h8d0;
      20'h046f2: out <= 12'h8d0;
      20'h046f3: out <= 12'h8d0;
      20'h046f4: out <= 12'h8d0;
      20'h046f5: out <= 12'h000;
      20'h046f6: out <= 12'h000;
      20'h046f7: out <= 12'h8d0;
      20'h046f8: out <= 12'h8d0;
      20'h046f9: out <= 12'h000;
      20'h046fa: out <= 12'h000;
      20'h046fb: out <= 12'h000;
      20'h046fc: out <= 12'h000;
      20'h046fd: out <= 12'h000;
      20'h046fe: out <= 12'h8d0;
      20'h046ff: out <= 12'h8d0;
      20'h04700: out <= 12'h8d0;
      20'h04701: out <= 12'h8d0;
      20'h04702: out <= 12'h000;
      20'h04703: out <= 12'h000;
      20'h04704: out <= 12'h8d0;
      20'h04705: out <= 12'h8d0;
      20'h04706: out <= 12'h000;
      20'h04707: out <= 12'h000;
      20'h04708: out <= 12'h000;
      20'h04709: out <= 12'h8d0;
      20'h0470a: out <= 12'h8d0;
      20'h0470b: out <= 12'h000;
      20'h0470c: out <= 12'h000;
      20'h0470d: out <= 12'h000;
      20'h0470e: out <= 12'h000;
      20'h0470f: out <= 12'h000;
      20'h04710: out <= 12'h000;
      20'h04711: out <= 12'h000;
      20'h04712: out <= 12'h000;
      20'h04713: out <= 12'h000;
      20'h04714: out <= 12'h000;
      20'h04715: out <= 12'h000;
      20'h04716: out <= 12'h000;
      20'h04717: out <= 12'h000;
      20'h04718: out <= 12'h603;
      20'h04719: out <= 12'h603;
      20'h0471a: out <= 12'h603;
      20'h0471b: out <= 12'h603;
      20'h0471c: out <= 12'h603;
      20'h0471d: out <= 12'h603;
      20'h0471e: out <= 12'h603;
      20'h0471f: out <= 12'h603;
      20'h04720: out <= 12'h603;
      20'h04721: out <= 12'h603;
      20'h04722: out <= 12'h603;
      20'h04723: out <= 12'h603;
      20'h04724: out <= 12'h603;
      20'h04725: out <= 12'h603;
      20'h04726: out <= 12'h603;
      20'h04727: out <= 12'h603;
      20'h04728: out <= 12'h603;
      20'h04729: out <= 12'h603;
      20'h0472a: out <= 12'h603;
      20'h0472b: out <= 12'h603;
      20'h0472c: out <= 12'h603;
      20'h0472d: out <= 12'h603;
      20'h0472e: out <= 12'h603;
      20'h0472f: out <= 12'h603;
      20'h04730: out <= 12'h603;
      20'h04731: out <= 12'h603;
      20'h04732: out <= 12'h603;
      20'h04733: out <= 12'h603;
      20'h04734: out <= 12'h603;
      20'h04735: out <= 12'h603;
      20'h04736: out <= 12'h603;
      20'h04737: out <= 12'h603;
      20'h04738: out <= 12'h603;
      20'h04739: out <= 12'h603;
      20'h0473a: out <= 12'h603;
      20'h0473b: out <= 12'h603;
      20'h0473c: out <= 12'h603;
      20'h0473d: out <= 12'h603;
      20'h0473e: out <= 12'h603;
      20'h0473f: out <= 12'h603;
      20'h04740: out <= 12'h603;
      20'h04741: out <= 12'h603;
      20'h04742: out <= 12'h603;
      20'h04743: out <= 12'h603;
      20'h04744: out <= 12'h603;
      20'h04745: out <= 12'h603;
      20'h04746: out <= 12'h603;
      20'h04747: out <= 12'h603;
      20'h04748: out <= 12'h603;
      20'h04749: out <= 12'h603;
      20'h0474a: out <= 12'h603;
      20'h0474b: out <= 12'h603;
      20'h0474c: out <= 12'h000;
      20'h0474d: out <= 12'h000;
      20'h0474e: out <= 12'h16d;
      20'h0474f: out <= 12'h6af;
      20'h04750: out <= 12'hfff;
      20'h04751: out <= 12'h6af;
      20'h04752: out <= 12'h16d;
      20'h04753: out <= 12'h000;
      20'h04754: out <= 12'h603;
      20'h04755: out <= 12'h603;
      20'h04756: out <= 12'h603;
      20'h04757: out <= 12'h603;
      20'h04758: out <= 12'h603;
      20'h04759: out <= 12'h603;
      20'h0475a: out <= 12'h603;
      20'h0475b: out <= 12'h603;
      20'h0475c: out <= 12'h603;
      20'h0475d: out <= 12'h603;
      20'h0475e: out <= 12'h603;
      20'h0475f: out <= 12'h603;
      20'h04760: out <= 12'h603;
      20'h04761: out <= 12'h603;
      20'h04762: out <= 12'h603;
      20'h04763: out <= 12'h603;
      20'h04764: out <= 12'h603;
      20'h04765: out <= 12'h603;
      20'h04766: out <= 12'h603;
      20'h04767: out <= 12'h603;
      20'h04768: out <= 12'h603;
      20'h04769: out <= 12'h603;
      20'h0476a: out <= 12'h603;
      20'h0476b: out <= 12'h603;
      20'h0476c: out <= 12'h000;
      20'h0476d: out <= 12'h000;
      20'h0476e: out <= 12'h660;
      20'h0476f: out <= 12'hbb0;
      20'h04770: out <= 12'hee9;
      20'h04771: out <= 12'hbb0;
      20'h04772: out <= 12'h660;
      20'h04773: out <= 12'h000;
      20'h04774: out <= 12'h603;
      20'h04775: out <= 12'h603;
      20'h04776: out <= 12'h603;
      20'h04777: out <= 12'h603;
      20'h04778: out <= 12'h222;
      20'h04779: out <= 12'h222;
      20'h0477a: out <= 12'h222;
      20'h0477b: out <= 12'h222;
      20'h0477c: out <= 12'h222;
      20'h0477d: out <= 12'h222;
      20'h0477e: out <= 12'h222;
      20'h0477f: out <= 12'h222;
      20'h04780: out <= 12'h222;
      20'h04781: out <= 12'h222;
      20'h04782: out <= 12'h222;
      20'h04783: out <= 12'h222;
      20'h04784: out <= 12'h222;
      20'h04785: out <= 12'h222;
      20'h04786: out <= 12'h222;
      20'h04787: out <= 12'h222;
      20'h04788: out <= 12'h000;
      20'h04789: out <= 12'h000;
      20'h0478a: out <= 12'h000;
      20'h0478b: out <= 12'h000;
      20'h0478c: out <= 12'h000;
      20'h0478d: out <= 12'h000;
      20'h0478e: out <= 12'h000;
      20'h0478f: out <= 12'h000;
      20'h04790: out <= 12'hbb0;
      20'h04791: out <= 12'h000;
      20'h04792: out <= 12'h000;
      20'h04793: out <= 12'h000;
      20'h04794: out <= 12'h000;
      20'h04795: out <= 12'h000;
      20'h04796: out <= 12'h000;
      20'h04797: out <= 12'h000;
      20'h04798: out <= 12'h603;
      20'h04799: out <= 12'h603;
      20'h0479a: out <= 12'h603;
      20'h0479b: out <= 12'h603;
      20'h0479c: out <= 12'h000;
      20'h0479d: out <= 12'h666;
      20'h0479e: out <= 12'hfff;
      20'h0479f: out <= 12'hfff;
      20'h047a0: out <= 12'hfff;
      20'h047a1: out <= 12'hfff;
      20'h047a2: out <= 12'hfff;
      20'h047a3: out <= 12'hfff;
      20'h047a4: out <= 12'hfff;
      20'h047a5: out <= 12'hfff;
      20'h047a6: out <= 12'hfff;
      20'h047a7: out <= 12'hfff;
      20'h047a8: out <= 12'hfff;
      20'h047a9: out <= 12'hfff;
      20'h047aa: out <= 12'hfff;
      20'h047ab: out <= 12'h666;
      20'h047ac: out <= 12'h000;
      20'h047ad: out <= 12'h000;
      20'h047ae: out <= 12'h000;
      20'h047af: out <= 12'hb27;
      20'h047b0: out <= 12'hb27;
      20'h047b1: out <= 12'hb27;
      20'h047b2: out <= 12'hb27;
      20'h047b3: out <= 12'hb27;
      20'h047b4: out <= 12'hb27;
      20'h047b5: out <= 12'hb27;
      20'h047b6: out <= 12'hb27;
      20'h047b7: out <= 12'hb27;
      20'h047b8: out <= 12'hb27;
      20'h047b9: out <= 12'hb27;
      20'h047ba: out <= 12'h000;
      20'h047bb: out <= 12'h000;
      20'h047bc: out <= 12'h000;
      20'h047bd: out <= 12'h000;
      20'h047be: out <= 12'h000;
      20'h047bf: out <= 12'h000;
      20'h047c0: out <= 12'h000;
      20'h047c1: out <= 12'h000;
      20'h047c2: out <= 12'h000;
      20'h047c3: out <= 12'hb27;
      20'h047c4: out <= 12'hb27;
      20'h047c5: out <= 12'hee9;
      20'h047c6: out <= 12'hee9;
      20'h047c7: out <= 12'h000;
      20'h047c8: out <= 12'h000;
      20'h047c9: out <= 12'h000;
      20'h047ca: out <= 12'h000;
      20'h047cb: out <= 12'h000;
      20'h047cc: out <= 12'h603;
      20'h047cd: out <= 12'h603;
      20'h047ce: out <= 12'h603;
      20'h047cf: out <= 12'h603;
      20'h047d0: out <= 12'h603;
      20'h047d1: out <= 12'h603;
      20'h047d2: out <= 12'h603;
      20'h047d3: out <= 12'h603;
      20'h047d4: out <= 12'h603;
      20'h047d5: out <= 12'h603;
      20'h047d6: out <= 12'h603;
      20'h047d7: out <= 12'h603;
      20'h047d8: out <= 12'h603;
      20'h047d9: out <= 12'h603;
      20'h047da: out <= 12'h603;
      20'h047db: out <= 12'h603;
      20'h047dc: out <= 12'h603;
      20'h047dd: out <= 12'h603;
      20'h047de: out <= 12'h603;
      20'h047df: out <= 12'h603;
      20'h047e0: out <= 12'h603;
      20'h047e1: out <= 12'h603;
      20'h047e2: out <= 12'h603;
      20'h047e3: out <= 12'h603;
      20'h047e4: out <= 12'h603;
      20'h047e5: out <= 12'h603;
      20'h047e6: out <= 12'h603;
      20'h047e7: out <= 12'h603;
      20'h047e8: out <= 12'h603;
      20'h047e9: out <= 12'h603;
      20'h047ea: out <= 12'h603;
      20'h047eb: out <= 12'h603;
      20'h047ec: out <= 12'h603;
      20'h047ed: out <= 12'h603;
      20'h047ee: out <= 12'h603;
      20'h047ef: out <= 12'h603;
      20'h047f0: out <= 12'hee9;
      20'h047f1: out <= 12'hf87;
      20'h047f2: out <= 12'hf87;
      20'h047f3: out <= 12'hf87;
      20'h047f4: out <= 12'hf87;
      20'h047f5: out <= 12'hf87;
      20'h047f6: out <= 12'hf87;
      20'h047f7: out <= 12'hb27;
      20'h047f8: out <= 12'h000;
      20'h047f9: out <= 12'h000;
      20'h047fa: out <= 12'h000;
      20'h047fb: out <= 12'h000;
      20'h047fc: out <= 12'h000;
      20'h047fd: out <= 12'h000;
      20'h047fe: out <= 12'h000;
      20'h047ff: out <= 12'h000;
      20'h04800: out <= 12'h000;
      20'h04801: out <= 12'h000;
      20'h04802: out <= 12'h8d0;
      20'h04803: out <= 12'h8d0;
      20'h04804: out <= 12'h8d0;
      20'h04805: out <= 12'h000;
      20'h04806: out <= 12'h000;
      20'h04807: out <= 12'h000;
      20'h04808: out <= 12'h8d0;
      20'h04809: out <= 12'h8d0;
      20'h0480a: out <= 12'h000;
      20'h0480b: out <= 12'h000;
      20'h0480c: out <= 12'h8d0;
      20'h0480d: out <= 12'h8d0;
      20'h0480e: out <= 12'h000;
      20'h0480f: out <= 12'h8d0;
      20'h04810: out <= 12'h8d0;
      20'h04811: out <= 12'h000;
      20'h04812: out <= 12'h000;
      20'h04813: out <= 12'h000;
      20'h04814: out <= 12'h000;
      20'h04815: out <= 12'h8d0;
      20'h04816: out <= 12'h8d0;
      20'h04817: out <= 12'h8d0;
      20'h04818: out <= 12'h8d0;
      20'h04819: out <= 12'h8d0;
      20'h0481a: out <= 12'h8d0;
      20'h0481b: out <= 12'h000;
      20'h0481c: out <= 12'h8d0;
      20'h0481d: out <= 12'h8d0;
      20'h0481e: out <= 12'h000;
      20'h0481f: out <= 12'h000;
      20'h04820: out <= 12'h000;
      20'h04821: out <= 12'h8d0;
      20'h04822: out <= 12'h8d0;
      20'h04823: out <= 12'h000;
      20'h04824: out <= 12'h000;
      20'h04825: out <= 12'h000;
      20'h04826: out <= 12'h000;
      20'h04827: out <= 12'h000;
      20'h04828: out <= 12'h000;
      20'h04829: out <= 12'h000;
      20'h0482a: out <= 12'h000;
      20'h0482b: out <= 12'h000;
      20'h0482c: out <= 12'h000;
      20'h0482d: out <= 12'h000;
      20'h0482e: out <= 12'h000;
      20'h0482f: out <= 12'h000;
      20'h04830: out <= 12'h603;
      20'h04831: out <= 12'h603;
      20'h04832: out <= 12'h603;
      20'h04833: out <= 12'h603;
      20'h04834: out <= 12'h603;
      20'h04835: out <= 12'h603;
      20'h04836: out <= 12'h603;
      20'h04837: out <= 12'h603;
      20'h04838: out <= 12'h603;
      20'h04839: out <= 12'h603;
      20'h0483a: out <= 12'h603;
      20'h0483b: out <= 12'h603;
      20'h0483c: out <= 12'h603;
      20'h0483d: out <= 12'h603;
      20'h0483e: out <= 12'h603;
      20'h0483f: out <= 12'h603;
      20'h04840: out <= 12'h603;
      20'h04841: out <= 12'h603;
      20'h04842: out <= 12'h603;
      20'h04843: out <= 12'h603;
      20'h04844: out <= 12'h603;
      20'h04845: out <= 12'h603;
      20'h04846: out <= 12'h603;
      20'h04847: out <= 12'h603;
      20'h04848: out <= 12'h603;
      20'h04849: out <= 12'h603;
      20'h0484a: out <= 12'h603;
      20'h0484b: out <= 12'h603;
      20'h0484c: out <= 12'h603;
      20'h0484d: out <= 12'h603;
      20'h0484e: out <= 12'h603;
      20'h0484f: out <= 12'h603;
      20'h04850: out <= 12'h603;
      20'h04851: out <= 12'h603;
      20'h04852: out <= 12'h603;
      20'h04853: out <= 12'h603;
      20'h04854: out <= 12'h603;
      20'h04855: out <= 12'h603;
      20'h04856: out <= 12'h603;
      20'h04857: out <= 12'h603;
      20'h04858: out <= 12'h603;
      20'h04859: out <= 12'h603;
      20'h0485a: out <= 12'h603;
      20'h0485b: out <= 12'h603;
      20'h0485c: out <= 12'h603;
      20'h0485d: out <= 12'h603;
      20'h0485e: out <= 12'h603;
      20'h0485f: out <= 12'h603;
      20'h04860: out <= 12'h603;
      20'h04861: out <= 12'h603;
      20'h04862: out <= 12'h603;
      20'h04863: out <= 12'h603;
      20'h04864: out <= 12'h000;
      20'h04865: out <= 12'h000;
      20'h04866: out <= 12'h16d;
      20'h04867: out <= 12'h6af;
      20'h04868: out <= 12'hfff;
      20'h04869: out <= 12'h6af;
      20'h0486a: out <= 12'h16d;
      20'h0486b: out <= 12'h000;
      20'h0486c: out <= 12'h603;
      20'h0486d: out <= 12'h603;
      20'h0486e: out <= 12'h603;
      20'h0486f: out <= 12'h603;
      20'h04870: out <= 12'h603;
      20'h04871: out <= 12'h603;
      20'h04872: out <= 12'h603;
      20'h04873: out <= 12'h603;
      20'h04874: out <= 12'h603;
      20'h04875: out <= 12'h603;
      20'h04876: out <= 12'h603;
      20'h04877: out <= 12'h603;
      20'h04878: out <= 12'h603;
      20'h04879: out <= 12'h603;
      20'h0487a: out <= 12'h603;
      20'h0487b: out <= 12'h603;
      20'h0487c: out <= 12'h603;
      20'h0487d: out <= 12'h603;
      20'h0487e: out <= 12'h603;
      20'h0487f: out <= 12'h603;
      20'h04880: out <= 12'h603;
      20'h04881: out <= 12'h603;
      20'h04882: out <= 12'h603;
      20'h04883: out <= 12'h603;
      20'h04884: out <= 12'h000;
      20'h04885: out <= 12'h000;
      20'h04886: out <= 12'h660;
      20'h04887: out <= 12'hbb0;
      20'h04888: out <= 12'hee9;
      20'h04889: out <= 12'hbb0;
      20'h0488a: out <= 12'h660;
      20'h0488b: out <= 12'h000;
      20'h0488c: out <= 12'h603;
      20'h0488d: out <= 12'h603;
      20'h0488e: out <= 12'h603;
      20'h0488f: out <= 12'h603;
      20'h04890: out <= 12'h222;
      20'h04891: out <= 12'h222;
      20'h04892: out <= 12'h222;
      20'h04893: out <= 12'h222;
      20'h04894: out <= 12'h222;
      20'h04895: out <= 12'h222;
      20'h04896: out <= 12'h222;
      20'h04897: out <= 12'h222;
      20'h04898: out <= 12'h222;
      20'h04899: out <= 12'h222;
      20'h0489a: out <= 12'h222;
      20'h0489b: out <= 12'h222;
      20'h0489c: out <= 12'h222;
      20'h0489d: out <= 12'h222;
      20'h0489e: out <= 12'h222;
      20'h0489f: out <= 12'h222;
      20'h048a0: out <= 12'h000;
      20'h048a1: out <= 12'h000;
      20'h048a2: out <= 12'h000;
      20'h048a3: out <= 12'h000;
      20'h048a4: out <= 12'h000;
      20'h048a5: out <= 12'h000;
      20'h048a6: out <= 12'h000;
      20'h048a7: out <= 12'h660;
      20'h048a8: out <= 12'hee9;
      20'h048a9: out <= 12'h660;
      20'h048aa: out <= 12'h000;
      20'h048ab: out <= 12'h000;
      20'h048ac: out <= 12'h000;
      20'h048ad: out <= 12'h000;
      20'h048ae: out <= 12'h000;
      20'h048af: out <= 12'h000;
      20'h048b0: out <= 12'h603;
      20'h048b1: out <= 12'h603;
      20'h048b2: out <= 12'h603;
      20'h048b3: out <= 12'h603;
      20'h048b4: out <= 12'h000;
      20'h048b5: out <= 12'h666;
      20'h048b6: out <= 12'hfff;
      20'h048b7: out <= 12'hfff;
      20'h048b8: out <= 12'h000;
      20'h048b9: out <= 12'hfff;
      20'h048ba: out <= 12'hfff;
      20'h048bb: out <= 12'h666;
      20'h048bc: out <= 12'h666;
      20'h048bd: out <= 12'h666;
      20'h048be: out <= 12'hfff;
      20'h048bf: out <= 12'hfff;
      20'h048c0: out <= 12'h000;
      20'h048c1: out <= 12'hfff;
      20'h048c2: out <= 12'hfff;
      20'h048c3: out <= 12'h666;
      20'h048c4: out <= 12'h000;
      20'h048c5: out <= 12'h000;
      20'h048c6: out <= 12'h000;
      20'h048c7: out <= 12'hb27;
      20'h048c8: out <= 12'hf87;
      20'h048c9: out <= 12'hee9;
      20'h048ca: out <= 12'hee9;
      20'h048cb: out <= 12'hf87;
      20'h048cc: out <= 12'hf87;
      20'h048cd: out <= 12'hf87;
      20'h048ce: out <= 12'hb27;
      20'h048cf: out <= 12'hb27;
      20'h048d0: out <= 12'hf87;
      20'h048d1: out <= 12'hee9;
      20'h048d2: out <= 12'h000;
      20'h048d3: out <= 12'h000;
      20'h048d4: out <= 12'h000;
      20'h048d5: out <= 12'h000;
      20'h048d6: out <= 12'h000;
      20'h048d7: out <= 12'h000;
      20'h048d8: out <= 12'h000;
      20'h048d9: out <= 12'h000;
      20'h048da: out <= 12'hb27;
      20'h048db: out <= 12'hf87;
      20'h048dc: out <= 12'hf87;
      20'h048dd: out <= 12'hb27;
      20'h048de: out <= 12'hb27;
      20'h048df: out <= 12'hee9;
      20'h048e0: out <= 12'hee9;
      20'h048e1: out <= 12'h000;
      20'h048e2: out <= 12'h000;
      20'h048e3: out <= 12'h000;
      20'h048e4: out <= 12'h603;
      20'h048e5: out <= 12'h603;
      20'h048e6: out <= 12'h603;
      20'h048e7: out <= 12'h603;
      20'h048e8: out <= 12'h603;
      20'h048e9: out <= 12'h603;
      20'h048ea: out <= 12'h603;
      20'h048eb: out <= 12'h603;
      20'h048ec: out <= 12'h603;
      20'h048ed: out <= 12'h603;
      20'h048ee: out <= 12'h603;
      20'h048ef: out <= 12'h603;
      20'h048f0: out <= 12'h603;
      20'h048f1: out <= 12'h603;
      20'h048f2: out <= 12'h603;
      20'h048f3: out <= 12'h603;
      20'h048f4: out <= 12'h603;
      20'h048f5: out <= 12'h603;
      20'h048f6: out <= 12'h603;
      20'h048f7: out <= 12'h603;
      20'h048f8: out <= 12'h603;
      20'h048f9: out <= 12'h603;
      20'h048fa: out <= 12'h603;
      20'h048fb: out <= 12'h603;
      20'h048fc: out <= 12'h603;
      20'h048fd: out <= 12'h603;
      20'h048fe: out <= 12'h603;
      20'h048ff: out <= 12'h603;
      20'h04900: out <= 12'h603;
      20'h04901: out <= 12'h603;
      20'h04902: out <= 12'h603;
      20'h04903: out <= 12'h603;
      20'h04904: out <= 12'h603;
      20'h04905: out <= 12'h603;
      20'h04906: out <= 12'h603;
      20'h04907: out <= 12'h603;
      20'h04908: out <= 12'hee9;
      20'h04909: out <= 12'hf87;
      20'h0490a: out <= 12'hee9;
      20'h0490b: out <= 12'hee9;
      20'h0490c: out <= 12'hee9;
      20'h0490d: out <= 12'hb27;
      20'h0490e: out <= 12'hf87;
      20'h0490f: out <= 12'hb27;
      20'h04910: out <= 12'h000;
      20'h04911: out <= 12'h000;
      20'h04912: out <= 12'h000;
      20'h04913: out <= 12'h000;
      20'h04914: out <= 12'h000;
      20'h04915: out <= 12'h000;
      20'h04916: out <= 12'h000;
      20'h04917: out <= 12'h000;
      20'h04918: out <= 12'h000;
      20'h04919: out <= 12'h000;
      20'h0491a: out <= 12'h000;
      20'h0491b: out <= 12'h8d0;
      20'h0491c: out <= 12'h8d0;
      20'h0491d: out <= 12'h000;
      20'h0491e: out <= 12'h000;
      20'h0491f: out <= 12'h000;
      20'h04920: out <= 12'h8d0;
      20'h04921: out <= 12'h8d0;
      20'h04922: out <= 12'h000;
      20'h04923: out <= 12'h000;
      20'h04924: out <= 12'h8d0;
      20'h04925: out <= 12'h8d0;
      20'h04926: out <= 12'h000;
      20'h04927: out <= 12'h8d0;
      20'h04928: out <= 12'h8d0;
      20'h04929: out <= 12'h000;
      20'h0492a: out <= 12'h000;
      20'h0492b: out <= 12'h000;
      20'h0492c: out <= 12'h000;
      20'h0492d: out <= 12'h8d0;
      20'h0492e: out <= 12'h8d0;
      20'h0492f: out <= 12'h000;
      20'h04930: out <= 12'h000;
      20'h04931: out <= 12'h8d0;
      20'h04932: out <= 12'h8d0;
      20'h04933: out <= 12'h000;
      20'h04934: out <= 12'h8d0;
      20'h04935: out <= 12'h8d0;
      20'h04936: out <= 12'h000;
      20'h04937: out <= 12'h000;
      20'h04938: out <= 12'h000;
      20'h04939: out <= 12'h8d0;
      20'h0493a: out <= 12'h8d0;
      20'h0493b: out <= 12'h000;
      20'h0493c: out <= 12'h000;
      20'h0493d: out <= 12'h000;
      20'h0493e: out <= 12'h000;
      20'h0493f: out <= 12'h000;
      20'h04940: out <= 12'h000;
      20'h04941: out <= 12'h000;
      20'h04942: out <= 12'h000;
      20'h04943: out <= 12'h000;
      20'h04944: out <= 12'h000;
      20'h04945: out <= 12'h000;
      20'h04946: out <= 12'h000;
      20'h04947: out <= 12'h000;
      20'h04948: out <= 12'h603;
      20'h04949: out <= 12'h603;
      20'h0494a: out <= 12'h603;
      20'h0494b: out <= 12'h603;
      20'h0494c: out <= 12'h603;
      20'h0494d: out <= 12'h603;
      20'h0494e: out <= 12'h603;
      20'h0494f: out <= 12'h603;
      20'h04950: out <= 12'h603;
      20'h04951: out <= 12'h603;
      20'h04952: out <= 12'h603;
      20'h04953: out <= 12'h603;
      20'h04954: out <= 12'h603;
      20'h04955: out <= 12'h603;
      20'h04956: out <= 12'h603;
      20'h04957: out <= 12'h603;
      20'h04958: out <= 12'h603;
      20'h04959: out <= 12'h603;
      20'h0495a: out <= 12'h603;
      20'h0495b: out <= 12'h603;
      20'h0495c: out <= 12'h603;
      20'h0495d: out <= 12'h603;
      20'h0495e: out <= 12'h603;
      20'h0495f: out <= 12'h603;
      20'h04960: out <= 12'h603;
      20'h04961: out <= 12'h603;
      20'h04962: out <= 12'h603;
      20'h04963: out <= 12'h603;
      20'h04964: out <= 12'h603;
      20'h04965: out <= 12'h603;
      20'h04966: out <= 12'h603;
      20'h04967: out <= 12'h603;
      20'h04968: out <= 12'h603;
      20'h04969: out <= 12'h603;
      20'h0496a: out <= 12'h603;
      20'h0496b: out <= 12'h603;
      20'h0496c: out <= 12'h603;
      20'h0496d: out <= 12'h603;
      20'h0496e: out <= 12'h603;
      20'h0496f: out <= 12'h603;
      20'h04970: out <= 12'h603;
      20'h04971: out <= 12'h603;
      20'h04972: out <= 12'h603;
      20'h04973: out <= 12'h603;
      20'h04974: out <= 12'h603;
      20'h04975: out <= 12'h603;
      20'h04976: out <= 12'h603;
      20'h04977: out <= 12'h603;
      20'h04978: out <= 12'h603;
      20'h04979: out <= 12'h603;
      20'h0497a: out <= 12'h603;
      20'h0497b: out <= 12'h603;
      20'h0497c: out <= 12'h000;
      20'h0497d: out <= 12'h000;
      20'h0497e: out <= 12'h16d;
      20'h0497f: out <= 12'h6af;
      20'h04980: out <= 12'hfff;
      20'h04981: out <= 12'h6af;
      20'h04982: out <= 12'h16d;
      20'h04983: out <= 12'h000;
      20'h04984: out <= 12'h603;
      20'h04985: out <= 12'h603;
      20'h04986: out <= 12'h603;
      20'h04987: out <= 12'h603;
      20'h04988: out <= 12'h603;
      20'h04989: out <= 12'h603;
      20'h0498a: out <= 12'h603;
      20'h0498b: out <= 12'h603;
      20'h0498c: out <= 12'h603;
      20'h0498d: out <= 12'h603;
      20'h0498e: out <= 12'h603;
      20'h0498f: out <= 12'h603;
      20'h04990: out <= 12'h603;
      20'h04991: out <= 12'h603;
      20'h04992: out <= 12'h603;
      20'h04993: out <= 12'h603;
      20'h04994: out <= 12'h603;
      20'h04995: out <= 12'h603;
      20'h04996: out <= 12'h603;
      20'h04997: out <= 12'h603;
      20'h04998: out <= 12'h603;
      20'h04999: out <= 12'h603;
      20'h0499a: out <= 12'h603;
      20'h0499b: out <= 12'h603;
      20'h0499c: out <= 12'h000;
      20'h0499d: out <= 12'h660;
      20'h0499e: out <= 12'hbb0;
      20'h0499f: out <= 12'hee9;
      20'h049a0: out <= 12'hee9;
      20'h049a1: out <= 12'hee9;
      20'h049a2: out <= 12'hbb0;
      20'h049a3: out <= 12'h660;
      20'h049a4: out <= 12'h603;
      20'h049a5: out <= 12'h603;
      20'h049a6: out <= 12'h603;
      20'h049a7: out <= 12'h603;
      20'h049a8: out <= 12'h222;
      20'h049a9: out <= 12'h222;
      20'h049aa: out <= 12'h222;
      20'h049ab: out <= 12'h222;
      20'h049ac: out <= 12'h660;
      20'h049ad: out <= 12'h222;
      20'h049ae: out <= 12'h222;
      20'h049af: out <= 12'h222;
      20'h049b0: out <= 12'h222;
      20'h049b1: out <= 12'h222;
      20'h049b2: out <= 12'h222;
      20'h049b3: out <= 12'h222;
      20'h049b4: out <= 12'h660;
      20'h049b5: out <= 12'h222;
      20'h049b6: out <= 12'h222;
      20'h049b7: out <= 12'h222;
      20'h049b8: out <= 12'h000;
      20'h049b9: out <= 12'h000;
      20'h049ba: out <= 12'h000;
      20'h049bb: out <= 12'h000;
      20'h049bc: out <= 12'h000;
      20'h049bd: out <= 12'h000;
      20'h049be: out <= 12'h660;
      20'h049bf: out <= 12'hbb0;
      20'h049c0: out <= 12'hee9;
      20'h049c1: out <= 12'hbb0;
      20'h049c2: out <= 12'h660;
      20'h049c3: out <= 12'h000;
      20'h049c4: out <= 12'h000;
      20'h049c5: out <= 12'h000;
      20'h049c6: out <= 12'h000;
      20'h049c7: out <= 12'h000;
      20'h049c8: out <= 12'h603;
      20'h049c9: out <= 12'h603;
      20'h049ca: out <= 12'h603;
      20'h049cb: out <= 12'h603;
      20'h049cc: out <= 12'h000;
      20'h049cd: out <= 12'h666;
      20'h049ce: out <= 12'hfff;
      20'h049cf: out <= 12'hfff;
      20'h049d0: out <= 12'hfff;
      20'h049d1: out <= 12'h000;
      20'h049d2: out <= 12'hfff;
      20'h049d3: out <= 12'hfff;
      20'h049d4: out <= 12'h666;
      20'h049d5: out <= 12'hfff;
      20'h049d6: out <= 12'hfff;
      20'h049d7: out <= 12'h000;
      20'h049d8: out <= 12'hfff;
      20'h049d9: out <= 12'hfff;
      20'h049da: out <= 12'hfff;
      20'h049db: out <= 12'h666;
      20'h049dc: out <= 12'h000;
      20'h049dd: out <= 12'h000;
      20'h049de: out <= 12'h000;
      20'h049df: out <= 12'hb27;
      20'h049e0: out <= 12'hf87;
      20'h049e1: out <= 12'hee9;
      20'h049e2: out <= 12'hee9;
      20'h049e3: out <= 12'hf87;
      20'h049e4: out <= 12'hf87;
      20'h049e5: out <= 12'hf87;
      20'h049e6: out <= 12'hb27;
      20'h049e7: out <= 12'hb27;
      20'h049e8: out <= 12'hf87;
      20'h049e9: out <= 12'hee9;
      20'h049ea: out <= 12'h000;
      20'h049eb: out <= 12'h000;
      20'h049ec: out <= 12'h000;
      20'h049ed: out <= 12'h000;
      20'h049ee: out <= 12'h000;
      20'h049ef: out <= 12'h000;
      20'h049f0: out <= 12'h000;
      20'h049f1: out <= 12'h000;
      20'h049f2: out <= 12'hb27;
      20'h049f3: out <= 12'hf87;
      20'h049f4: out <= 12'hee9;
      20'h049f5: out <= 12'hee9;
      20'h049f6: out <= 12'hf87;
      20'h049f7: out <= 12'hb27;
      20'h049f8: out <= 12'hb27;
      20'h049f9: out <= 12'hee9;
      20'h049fa: out <= 12'hee9;
      20'h049fb: out <= 12'h000;
      20'h049fc: out <= 12'h603;
      20'h049fd: out <= 12'h603;
      20'h049fe: out <= 12'h603;
      20'h049ff: out <= 12'h603;
      20'h04a00: out <= 12'h603;
      20'h04a01: out <= 12'h603;
      20'h04a02: out <= 12'h603;
      20'h04a03: out <= 12'h603;
      20'h04a04: out <= 12'h603;
      20'h04a05: out <= 12'h603;
      20'h04a06: out <= 12'h603;
      20'h04a07: out <= 12'h603;
      20'h04a08: out <= 12'h603;
      20'h04a09: out <= 12'h603;
      20'h04a0a: out <= 12'h603;
      20'h04a0b: out <= 12'h603;
      20'h04a0c: out <= 12'h603;
      20'h04a0d: out <= 12'h603;
      20'h04a0e: out <= 12'h603;
      20'h04a0f: out <= 12'h603;
      20'h04a10: out <= 12'h603;
      20'h04a11: out <= 12'h603;
      20'h04a12: out <= 12'h603;
      20'h04a13: out <= 12'h603;
      20'h04a14: out <= 12'h603;
      20'h04a15: out <= 12'h603;
      20'h04a16: out <= 12'h603;
      20'h04a17: out <= 12'h603;
      20'h04a18: out <= 12'h603;
      20'h04a19: out <= 12'h603;
      20'h04a1a: out <= 12'h603;
      20'h04a1b: out <= 12'h603;
      20'h04a1c: out <= 12'h603;
      20'h04a1d: out <= 12'h603;
      20'h04a1e: out <= 12'h603;
      20'h04a1f: out <= 12'h603;
      20'h04a20: out <= 12'hee9;
      20'h04a21: out <= 12'hf87;
      20'h04a22: out <= 12'hee9;
      20'h04a23: out <= 12'hf87;
      20'h04a24: out <= 12'hf87;
      20'h04a25: out <= 12'hb27;
      20'h04a26: out <= 12'hf87;
      20'h04a27: out <= 12'hb27;
      20'h04a28: out <= 12'h000;
      20'h04a29: out <= 12'h000;
      20'h04a2a: out <= 12'h000;
      20'h04a2b: out <= 12'h000;
      20'h04a2c: out <= 12'h000;
      20'h04a2d: out <= 12'h000;
      20'h04a2e: out <= 12'h000;
      20'h04a2f: out <= 12'h000;
      20'h04a30: out <= 12'h000;
      20'h04a31: out <= 12'h000;
      20'h04a32: out <= 12'h000;
      20'h04a33: out <= 12'h8d0;
      20'h04a34: out <= 12'h8d0;
      20'h04a35: out <= 12'h000;
      20'h04a36: out <= 12'h000;
      20'h04a37: out <= 12'h000;
      20'h04a38: out <= 12'h8d0;
      20'h04a39: out <= 12'h8d0;
      20'h04a3a: out <= 12'h8d0;
      20'h04a3b: out <= 12'h8d0;
      20'h04a3c: out <= 12'h8d0;
      20'h04a3d: out <= 12'h000;
      20'h04a3e: out <= 12'h000;
      20'h04a3f: out <= 12'h8d0;
      20'h04a40: out <= 12'h8d0;
      20'h04a41: out <= 12'h000;
      20'h04a42: out <= 12'h000;
      20'h04a43: out <= 12'h000;
      20'h04a44: out <= 12'h000;
      20'h04a45: out <= 12'h8d0;
      20'h04a46: out <= 12'h8d0;
      20'h04a47: out <= 12'h000;
      20'h04a48: out <= 12'h000;
      20'h04a49: out <= 12'h8d0;
      20'h04a4a: out <= 12'h8d0;
      20'h04a4b: out <= 12'h000;
      20'h04a4c: out <= 12'h000;
      20'h04a4d: out <= 12'h8d0;
      20'h04a4e: out <= 12'h8d0;
      20'h04a4f: out <= 12'h8d0;
      20'h04a50: out <= 12'h8d0;
      20'h04a51: out <= 12'h8d0;
      20'h04a52: out <= 12'h000;
      20'h04a53: out <= 12'h000;
      20'h04a54: out <= 12'h000;
      20'h04a55: out <= 12'h000;
      20'h04a56: out <= 12'h000;
      20'h04a57: out <= 12'h000;
      20'h04a58: out <= 12'h000;
      20'h04a59: out <= 12'h000;
      20'h04a5a: out <= 12'h000;
      20'h04a5b: out <= 12'h000;
      20'h04a5c: out <= 12'h000;
      20'h04a5d: out <= 12'h000;
      20'h04a5e: out <= 12'h000;
      20'h04a5f: out <= 12'h000;
      20'h04a60: out <= 12'h603;
      20'h04a61: out <= 12'h603;
      20'h04a62: out <= 12'h603;
      20'h04a63: out <= 12'h603;
      20'h04a64: out <= 12'h222;
      20'h04a65: out <= 12'h222;
      20'h04a66: out <= 12'h222;
      20'h04a67: out <= 12'h222;
      20'h04a68: out <= 12'h222;
      20'h04a69: out <= 12'h222;
      20'h04a6a: out <= 12'h222;
      20'h04a6b: out <= 12'h222;
      20'h04a6c: out <= 12'h603;
      20'h04a6d: out <= 12'h603;
      20'h04a6e: out <= 12'h603;
      20'h04a6f: out <= 12'h603;
      20'h04a70: out <= 12'h603;
      20'h04a71: out <= 12'h603;
      20'h04a72: out <= 12'h603;
      20'h04a73: out <= 12'h603;
      20'h04a74: out <= 12'h000;
      20'h04a75: out <= 12'h000;
      20'h04a76: out <= 12'h000;
      20'h04a77: out <= 12'h6af;
      20'h04a78: out <= 12'h6af;
      20'h04a79: out <= 12'h000;
      20'h04a7a: out <= 12'h000;
      20'h04a7b: out <= 12'h000;
      20'h04a7c: out <= 12'h603;
      20'h04a7d: out <= 12'h603;
      20'h04a7e: out <= 12'h603;
      20'h04a7f: out <= 12'h603;
      20'h04a80: out <= 12'h222;
      20'h04a81: out <= 12'h6af;
      20'h04a82: out <= 12'h6af;
      20'h04a83: out <= 12'h222;
      20'h04a84: out <= 12'h222;
      20'h04a85: out <= 12'h222;
      20'h04a86: out <= 12'h222;
      20'h04a87: out <= 12'h222;
      20'h04a88: out <= 12'h222;
      20'h04a89: out <= 12'h222;
      20'h04a8a: out <= 12'h222;
      20'h04a8b: out <= 12'h222;
      20'h04a8c: out <= 12'h222;
      20'h04a8d: out <= 12'h222;
      20'h04a8e: out <= 12'h222;
      20'h04a8f: out <= 12'h222;
      20'h04a90: out <= 12'h603;
      20'h04a91: out <= 12'h603;
      20'h04a92: out <= 12'h603;
      20'h04a93: out <= 12'h603;
      20'h04a94: out <= 12'h000;
      20'h04a95: out <= 12'h000;
      20'h04a96: out <= 12'h16d;
      20'h04a97: out <= 12'h6af;
      20'h04a98: out <= 12'hfff;
      20'h04a99: out <= 12'h6af;
      20'h04a9a: out <= 12'h16d;
      20'h04a9b: out <= 12'h000;
      20'h04a9c: out <= 12'h603;
      20'h04a9d: out <= 12'h603;
      20'h04a9e: out <= 12'h603;
      20'h04a9f: out <= 12'h603;
      20'h04aa0: out <= 12'h222;
      20'h04aa1: out <= 12'h222;
      20'h04aa2: out <= 12'h222;
      20'h04aa3: out <= 12'h222;
      20'h04aa4: out <= 12'h222;
      20'h04aa5: out <= 12'h222;
      20'h04aa6: out <= 12'h222;
      20'h04aa7: out <= 12'h222;
      20'h04aa8: out <= 12'h660;
      20'h04aa9: out <= 12'h660;
      20'h04aaa: out <= 12'h660;
      20'h04aab: out <= 12'h660;
      20'h04aac: out <= 12'h660;
      20'h04aad: out <= 12'h222;
      20'h04aae: out <= 12'h222;
      20'h04aaf: out <= 12'h222;
      20'h04ab0: out <= 12'h603;
      20'h04ab1: out <= 12'h603;
      20'h04ab2: out <= 12'h603;
      20'h04ab3: out <= 12'h603;
      20'h04ab4: out <= 12'h000;
      20'h04ab5: out <= 12'h660;
      20'h04ab6: out <= 12'hbb0;
      20'h04ab7: out <= 12'hee9;
      20'h04ab8: out <= 12'hee9;
      20'h04ab9: out <= 12'hee9;
      20'h04aba: out <= 12'hbb0;
      20'h04abb: out <= 12'h660;
      20'h04abc: out <= 12'h603;
      20'h04abd: out <= 12'h603;
      20'h04abe: out <= 12'h603;
      20'h04abf: out <= 12'h603;
      20'h04ac0: out <= 12'h222;
      20'h04ac1: out <= 12'h222;
      20'h04ac2: out <= 12'h222;
      20'h04ac3: out <= 12'h222;
      20'h04ac4: out <= 12'h222;
      20'h04ac5: out <= 12'hbb0;
      20'h04ac6: out <= 12'h222;
      20'h04ac7: out <= 12'h660;
      20'h04ac8: out <= 12'h660;
      20'h04ac9: out <= 12'h660;
      20'h04aca: out <= 12'h222;
      20'h04acb: out <= 12'hbb0;
      20'h04acc: out <= 12'h222;
      20'h04acd: out <= 12'h222;
      20'h04ace: out <= 12'h222;
      20'h04acf: out <= 12'h222;
      20'h04ad0: out <= 12'h000;
      20'h04ad1: out <= 12'h000;
      20'h04ad2: out <= 12'h000;
      20'h04ad3: out <= 12'h000;
      20'h04ad4: out <= 12'h000;
      20'h04ad5: out <= 12'h660;
      20'h04ad6: out <= 12'hbb0;
      20'h04ad7: out <= 12'hee9;
      20'h04ad8: out <= 12'hee9;
      20'h04ad9: out <= 12'hee9;
      20'h04ada: out <= 12'hbb0;
      20'h04adb: out <= 12'h660;
      20'h04adc: out <= 12'h000;
      20'h04add: out <= 12'h000;
      20'h04ade: out <= 12'h000;
      20'h04adf: out <= 12'h000;
      20'h04ae0: out <= 12'h603;
      20'h04ae1: out <= 12'h603;
      20'h04ae2: out <= 12'h603;
      20'h04ae3: out <= 12'h603;
      20'h04ae4: out <= 12'h000;
      20'h04ae5: out <= 12'h666;
      20'h04ae6: out <= 12'hfff;
      20'h04ae7: out <= 12'h666;
      20'h04ae8: out <= 12'h666;
      20'h04ae9: out <= 12'hfff;
      20'h04aea: out <= 12'h000;
      20'h04aeb: out <= 12'hfff;
      20'h04aec: out <= 12'h666;
      20'h04aed: out <= 12'hfff;
      20'h04aee: out <= 12'h000;
      20'h04aef: out <= 12'hfff;
      20'h04af0: out <= 12'h666;
      20'h04af1: out <= 12'h666;
      20'h04af2: out <= 12'hfff;
      20'h04af3: out <= 12'h666;
      20'h04af4: out <= 12'h000;
      20'h04af5: out <= 12'h000;
      20'h04af6: out <= 12'h000;
      20'h04af7: out <= 12'hb27;
      20'h04af8: out <= 12'hf87;
      20'h04af9: out <= 12'hee9;
      20'h04afa: out <= 12'hee9;
      20'h04afb: out <= 12'hf87;
      20'h04afc: out <= 12'hf87;
      20'h04afd: out <= 12'hf87;
      20'h04afe: out <= 12'hb27;
      20'h04aff: out <= 12'hb27;
      20'h04b00: out <= 12'hf87;
      20'h04b01: out <= 12'hee9;
      20'h04b02: out <= 12'h000;
      20'h04b03: out <= 12'h000;
      20'h04b04: out <= 12'h000;
      20'h04b05: out <= 12'h000;
      20'h04b06: out <= 12'h000;
      20'h04b07: out <= 12'h000;
      20'h04b08: out <= 12'h000;
      20'h04b09: out <= 12'hb27;
      20'h04b0a: out <= 12'hf87;
      20'h04b0b: out <= 12'hee9;
      20'h04b0c: out <= 12'hee9;
      20'h04b0d: out <= 12'hf87;
      20'h04b0e: out <= 12'hf87;
      20'h04b0f: out <= 12'hf87;
      20'h04b10: out <= 12'hb27;
      20'h04b11: out <= 12'hb27;
      20'h04b12: out <= 12'hb27;
      20'h04b13: out <= 12'hee9;
      20'h04b14: out <= 12'h603;
      20'h04b15: out <= 12'h603;
      20'h04b16: out <= 12'h603;
      20'h04b17: out <= 12'h603;
      20'h04b18: out <= 12'h603;
      20'h04b19: out <= 12'h603;
      20'h04b1a: out <= 12'h603;
      20'h04b1b: out <= 12'h603;
      20'h04b1c: out <= 12'h603;
      20'h04b1d: out <= 12'h603;
      20'h04b1e: out <= 12'h603;
      20'h04b1f: out <= 12'h603;
      20'h04b20: out <= 12'h603;
      20'h04b21: out <= 12'h603;
      20'h04b22: out <= 12'h603;
      20'h04b23: out <= 12'h603;
      20'h04b24: out <= 12'h603;
      20'h04b25: out <= 12'h603;
      20'h04b26: out <= 12'h603;
      20'h04b27: out <= 12'h603;
      20'h04b28: out <= 12'h603;
      20'h04b29: out <= 12'h603;
      20'h04b2a: out <= 12'h603;
      20'h04b2b: out <= 12'h603;
      20'h04b2c: out <= 12'h603;
      20'h04b2d: out <= 12'h603;
      20'h04b2e: out <= 12'h603;
      20'h04b2f: out <= 12'h603;
      20'h04b30: out <= 12'h603;
      20'h04b31: out <= 12'h603;
      20'h04b32: out <= 12'h603;
      20'h04b33: out <= 12'h603;
      20'h04b34: out <= 12'h603;
      20'h04b35: out <= 12'h603;
      20'h04b36: out <= 12'h603;
      20'h04b37: out <= 12'h603;
      20'h04b38: out <= 12'hee9;
      20'h04b39: out <= 12'hf87;
      20'h04b3a: out <= 12'hee9;
      20'h04b3b: out <= 12'hf87;
      20'h04b3c: out <= 12'hf87;
      20'h04b3d: out <= 12'hb27;
      20'h04b3e: out <= 12'hf87;
      20'h04b3f: out <= 12'hb27;
      20'h04b40: out <= 12'h000;
      20'h04b41: out <= 12'h000;
      20'h04b42: out <= 12'h000;
      20'h04b43: out <= 12'h000;
      20'h04b44: out <= 12'h000;
      20'h04b45: out <= 12'h000;
      20'h04b46: out <= 12'h000;
      20'h04b47: out <= 12'h000;
      20'h04b48: out <= 12'h000;
      20'h04b49: out <= 12'h000;
      20'h04b4a: out <= 12'h000;
      20'h04b4b: out <= 12'h8d0;
      20'h04b4c: out <= 12'h8d0;
      20'h04b4d: out <= 12'h000;
      20'h04b4e: out <= 12'h000;
      20'h04b4f: out <= 12'h000;
      20'h04b50: out <= 12'h8d0;
      20'h04b51: out <= 12'h8d0;
      20'h04b52: out <= 12'h000;
      20'h04b53: out <= 12'h000;
      20'h04b54: out <= 12'h000;
      20'h04b55: out <= 12'h000;
      20'h04b56: out <= 12'h000;
      20'h04b57: out <= 12'h8d0;
      20'h04b58: out <= 12'h8d0;
      20'h04b59: out <= 12'h000;
      20'h04b5a: out <= 12'h000;
      20'h04b5b: out <= 12'h000;
      20'h04b5c: out <= 12'h000;
      20'h04b5d: out <= 12'h8d0;
      20'h04b5e: out <= 12'h8d0;
      20'h04b5f: out <= 12'h8d0;
      20'h04b60: out <= 12'h8d0;
      20'h04b61: out <= 12'h8d0;
      20'h04b62: out <= 12'h8d0;
      20'h04b63: out <= 12'h000;
      20'h04b64: out <= 12'h000;
      20'h04b65: out <= 12'h000;
      20'h04b66: out <= 12'h8d0;
      20'h04b67: out <= 12'h8d0;
      20'h04b68: out <= 12'h8d0;
      20'h04b69: out <= 12'h000;
      20'h04b6a: out <= 12'h000;
      20'h04b6b: out <= 12'h000;
      20'h04b6c: out <= 12'h000;
      20'h04b6d: out <= 12'h000;
      20'h04b6e: out <= 12'h000;
      20'h04b6f: out <= 12'h000;
      20'h04b70: out <= 12'h000;
      20'h04b71: out <= 12'h000;
      20'h04b72: out <= 12'h000;
      20'h04b73: out <= 12'h000;
      20'h04b74: out <= 12'h000;
      20'h04b75: out <= 12'h000;
      20'h04b76: out <= 12'h000;
      20'h04b77: out <= 12'h000;
      20'h04b78: out <= 12'h603;
      20'h04b79: out <= 12'h603;
      20'h04b7a: out <= 12'h603;
      20'h04b7b: out <= 12'h603;
      20'h04b7c: out <= 12'h222;
      20'h04b7d: out <= 12'h222;
      20'h04b7e: out <= 12'h222;
      20'h04b7f: out <= 12'h222;
      20'h04b80: out <= 12'h222;
      20'h04b81: out <= 12'h222;
      20'h04b82: out <= 12'h222;
      20'h04b83: out <= 12'h222;
      20'h04b84: out <= 12'h603;
      20'h04b85: out <= 12'h603;
      20'h04b86: out <= 12'h603;
      20'h04b87: out <= 12'h603;
      20'h04b88: out <= 12'h603;
      20'h04b89: out <= 12'h603;
      20'h04b8a: out <= 12'h603;
      20'h04b8b: out <= 12'h603;
      20'h04b8c: out <= 12'h000;
      20'h04b8d: out <= 12'h000;
      20'h04b8e: out <= 12'h000;
      20'h04b8f: out <= 12'h6af;
      20'h04b90: out <= 12'h6af;
      20'h04b91: out <= 12'h000;
      20'h04b92: out <= 12'h000;
      20'h04b93: out <= 12'h000;
      20'h04b94: out <= 12'h603;
      20'h04b95: out <= 12'h603;
      20'h04b96: out <= 12'h603;
      20'h04b97: out <= 12'h603;
      20'h04b98: out <= 12'h222;
      20'h04b99: out <= 12'h16d;
      20'h04b9a: out <= 12'h16d;
      20'h04b9b: out <= 12'h16d;
      20'h04b9c: out <= 12'h222;
      20'h04b9d: out <= 12'h16d;
      20'h04b9e: out <= 12'h16d;
      20'h04b9f: out <= 12'h16d;
      20'h04ba0: out <= 12'h16d;
      20'h04ba1: out <= 12'h16d;
      20'h04ba2: out <= 12'h16d;
      20'h04ba3: out <= 12'h16d;
      20'h04ba4: out <= 12'h16d;
      20'h04ba5: out <= 12'h16d;
      20'h04ba6: out <= 12'h16d;
      20'h04ba7: out <= 12'h222;
      20'h04ba8: out <= 12'h603;
      20'h04ba9: out <= 12'h603;
      20'h04baa: out <= 12'h603;
      20'h04bab: out <= 12'h603;
      20'h04bac: out <= 12'h000;
      20'h04bad: out <= 12'h000;
      20'h04bae: out <= 12'h16d;
      20'h04baf: out <= 12'h6af;
      20'h04bb0: out <= 12'hfff;
      20'h04bb1: out <= 12'h6af;
      20'h04bb2: out <= 12'h16d;
      20'h04bb3: out <= 12'h000;
      20'h04bb4: out <= 12'h603;
      20'h04bb5: out <= 12'h603;
      20'h04bb6: out <= 12'h603;
      20'h04bb7: out <= 12'h603;
      20'h04bb8: out <= 12'h222;
      20'h04bb9: out <= 12'h222;
      20'h04bba: out <= 12'h222;
      20'h04bbb: out <= 12'h222;
      20'h04bbc: out <= 12'h222;
      20'h04bbd: out <= 12'h222;
      20'h04bbe: out <= 12'h660;
      20'h04bbf: out <= 12'h660;
      20'h04bc0: out <= 12'hbb0;
      20'h04bc1: out <= 12'hbb0;
      20'h04bc2: out <= 12'hbb0;
      20'h04bc3: out <= 12'hbb0;
      20'h04bc4: out <= 12'hbb0;
      20'h04bc5: out <= 12'h660;
      20'h04bc6: out <= 12'h660;
      20'h04bc7: out <= 12'h222;
      20'h04bc8: out <= 12'h603;
      20'h04bc9: out <= 12'h603;
      20'h04bca: out <= 12'h603;
      20'h04bcb: out <= 12'h603;
      20'h04bcc: out <= 12'h000;
      20'h04bcd: out <= 12'h660;
      20'h04bce: out <= 12'hbb0;
      20'h04bcf: out <= 12'hee9;
      20'h04bd0: out <= 12'hee9;
      20'h04bd1: out <= 12'hee9;
      20'h04bd2: out <= 12'hbb0;
      20'h04bd3: out <= 12'h660;
      20'h04bd4: out <= 12'h603;
      20'h04bd5: out <= 12'h603;
      20'h04bd6: out <= 12'h603;
      20'h04bd7: out <= 12'h603;
      20'h04bd8: out <= 12'h222;
      20'h04bd9: out <= 12'h222;
      20'h04bda: out <= 12'h222;
      20'h04bdb: out <= 12'h222;
      20'h04bdc: out <= 12'h222;
      20'h04bdd: out <= 12'h222;
      20'h04bde: out <= 12'hee9;
      20'h04bdf: out <= 12'hbb0;
      20'h04be0: out <= 12'hbb0;
      20'h04be1: out <= 12'hbb0;
      20'h04be2: out <= 12'hee9;
      20'h04be3: out <= 12'h222;
      20'h04be4: out <= 12'h222;
      20'h04be5: out <= 12'h222;
      20'h04be6: out <= 12'h222;
      20'h04be7: out <= 12'h222;
      20'h04be8: out <= 12'h000;
      20'h04be9: out <= 12'h000;
      20'h04bea: out <= 12'h000;
      20'h04beb: out <= 12'h000;
      20'h04bec: out <= 12'h660;
      20'h04bed: out <= 12'hbb0;
      20'h04bee: out <= 12'hee9;
      20'h04bef: out <= 12'hee9;
      20'h04bf0: out <= 12'hee9;
      20'h04bf1: out <= 12'hee9;
      20'h04bf2: out <= 12'hee9;
      20'h04bf3: out <= 12'hbb0;
      20'h04bf4: out <= 12'h660;
      20'h04bf5: out <= 12'h000;
      20'h04bf6: out <= 12'h000;
      20'h04bf7: out <= 12'h000;
      20'h04bf8: out <= 12'h603;
      20'h04bf9: out <= 12'h603;
      20'h04bfa: out <= 12'h603;
      20'h04bfb: out <= 12'h603;
      20'h04bfc: out <= 12'h000;
      20'h04bfd: out <= 12'h666;
      20'h04bfe: out <= 12'hfff;
      20'h04bff: out <= 12'h666;
      20'h04c00: out <= 12'h666;
      20'h04c01: out <= 12'hfff;
      20'h04c02: out <= 12'h666;
      20'h04c03: out <= 12'h000;
      20'h04c04: out <= 12'h666;
      20'h04c05: out <= 12'h000;
      20'h04c06: out <= 12'h666;
      20'h04c07: out <= 12'hfff;
      20'h04c08: out <= 12'h666;
      20'h04c09: out <= 12'h666;
      20'h04c0a: out <= 12'hfff;
      20'h04c0b: out <= 12'h666;
      20'h04c0c: out <= 12'h000;
      20'h04c0d: out <= 12'h000;
      20'h04c0e: out <= 12'h000;
      20'h04c0f: out <= 12'hb27;
      20'h04c10: out <= 12'hf87;
      20'h04c11: out <= 12'hee9;
      20'h04c12: out <= 12'hee9;
      20'h04c13: out <= 12'hf87;
      20'h04c14: out <= 12'hf87;
      20'h04c15: out <= 12'hf87;
      20'h04c16: out <= 12'hb27;
      20'h04c17: out <= 12'hb27;
      20'h04c18: out <= 12'hf87;
      20'h04c19: out <= 12'hee9;
      20'h04c1a: out <= 12'h000;
      20'h04c1b: out <= 12'h000;
      20'h04c1c: out <= 12'h000;
      20'h04c1d: out <= 12'h000;
      20'h04c1e: out <= 12'h000;
      20'h04c1f: out <= 12'h000;
      20'h04c20: out <= 12'h000;
      20'h04c21: out <= 12'hb27;
      20'h04c22: out <= 12'hf87;
      20'h04c23: out <= 12'hee9;
      20'h04c24: out <= 12'hee9;
      20'h04c25: out <= 12'hf87;
      20'h04c26: out <= 12'hf87;
      20'h04c27: out <= 12'hb27;
      20'h04c28: out <= 12'hb27;
      20'h04c29: out <= 12'hb27;
      20'h04c2a: out <= 12'hf87;
      20'h04c2b: out <= 12'h000;
      20'h04c2c: out <= 12'h603;
      20'h04c2d: out <= 12'h603;
      20'h04c2e: out <= 12'h603;
      20'h04c2f: out <= 12'h603;
      20'h04c30: out <= 12'h603;
      20'h04c31: out <= 12'h603;
      20'h04c32: out <= 12'h603;
      20'h04c33: out <= 12'h603;
      20'h04c34: out <= 12'h603;
      20'h04c35: out <= 12'h603;
      20'h04c36: out <= 12'h603;
      20'h04c37: out <= 12'h603;
      20'h04c38: out <= 12'h603;
      20'h04c39: out <= 12'h603;
      20'h04c3a: out <= 12'h603;
      20'h04c3b: out <= 12'h603;
      20'h04c3c: out <= 12'h603;
      20'h04c3d: out <= 12'h603;
      20'h04c3e: out <= 12'h603;
      20'h04c3f: out <= 12'h603;
      20'h04c40: out <= 12'h603;
      20'h04c41: out <= 12'h603;
      20'h04c42: out <= 12'h603;
      20'h04c43: out <= 12'h603;
      20'h04c44: out <= 12'h603;
      20'h04c45: out <= 12'h603;
      20'h04c46: out <= 12'h603;
      20'h04c47: out <= 12'h603;
      20'h04c48: out <= 12'h603;
      20'h04c49: out <= 12'h603;
      20'h04c4a: out <= 12'h603;
      20'h04c4b: out <= 12'h603;
      20'h04c4c: out <= 12'h603;
      20'h04c4d: out <= 12'h603;
      20'h04c4e: out <= 12'h603;
      20'h04c4f: out <= 12'h603;
      20'h04c50: out <= 12'hee9;
      20'h04c51: out <= 12'hf87;
      20'h04c52: out <= 12'hee9;
      20'h04c53: out <= 12'hb27;
      20'h04c54: out <= 12'hb27;
      20'h04c55: out <= 12'hb27;
      20'h04c56: out <= 12'hf87;
      20'h04c57: out <= 12'hb27;
      20'h04c58: out <= 12'h000;
      20'h04c59: out <= 12'h000;
      20'h04c5a: out <= 12'h000;
      20'h04c5b: out <= 12'h000;
      20'h04c5c: out <= 12'h000;
      20'h04c5d: out <= 12'h000;
      20'h04c5e: out <= 12'h000;
      20'h04c5f: out <= 12'h000;
      20'h04c60: out <= 12'h000;
      20'h04c61: out <= 12'h000;
      20'h04c62: out <= 12'h000;
      20'h04c63: out <= 12'h8d0;
      20'h04c64: out <= 12'h8d0;
      20'h04c65: out <= 12'h000;
      20'h04c66: out <= 12'h000;
      20'h04c67: out <= 12'h000;
      20'h04c68: out <= 12'h8d0;
      20'h04c69: out <= 12'h8d0;
      20'h04c6a: out <= 12'h000;
      20'h04c6b: out <= 12'h000;
      20'h04c6c: out <= 12'h000;
      20'h04c6d: out <= 12'h000;
      20'h04c6e: out <= 12'h000;
      20'h04c6f: out <= 12'h8d0;
      20'h04c70: out <= 12'h8d0;
      20'h04c71: out <= 12'h000;
      20'h04c72: out <= 12'h000;
      20'h04c73: out <= 12'h000;
      20'h04c74: out <= 12'h000;
      20'h04c75: out <= 12'h8d0;
      20'h04c76: out <= 12'h8d0;
      20'h04c77: out <= 12'h000;
      20'h04c78: out <= 12'h000;
      20'h04c79: out <= 12'h8d0;
      20'h04c7a: out <= 12'h8d0;
      20'h04c7b: out <= 12'h000;
      20'h04c7c: out <= 12'h000;
      20'h04c7d: out <= 12'h000;
      20'h04c7e: out <= 12'h8d0;
      20'h04c7f: out <= 12'h8d0;
      20'h04c80: out <= 12'h8d0;
      20'h04c81: out <= 12'h000;
      20'h04c82: out <= 12'h000;
      20'h04c83: out <= 12'h000;
      20'h04c84: out <= 12'h000;
      20'h04c85: out <= 12'h000;
      20'h04c86: out <= 12'h000;
      20'h04c87: out <= 12'h000;
      20'h04c88: out <= 12'h000;
      20'h04c89: out <= 12'h000;
      20'h04c8a: out <= 12'h000;
      20'h04c8b: out <= 12'h000;
      20'h04c8c: out <= 12'h000;
      20'h04c8d: out <= 12'h000;
      20'h04c8e: out <= 12'h000;
      20'h04c8f: out <= 12'h000;
      20'h04c90: out <= 12'h603;
      20'h04c91: out <= 12'h603;
      20'h04c92: out <= 12'h603;
      20'h04c93: out <= 12'h603;
      20'h04c94: out <= 12'h222;
      20'h04c95: out <= 12'h222;
      20'h04c96: out <= 12'h222;
      20'h04c97: out <= 12'h222;
      20'h04c98: out <= 12'h222;
      20'h04c99: out <= 12'h222;
      20'h04c9a: out <= 12'h222;
      20'h04c9b: out <= 12'h222;
      20'h04c9c: out <= 12'h603;
      20'h04c9d: out <= 12'h603;
      20'h04c9e: out <= 12'h603;
      20'h04c9f: out <= 12'h603;
      20'h04ca0: out <= 12'h603;
      20'h04ca1: out <= 12'h603;
      20'h04ca2: out <= 12'h603;
      20'h04ca3: out <= 12'h603;
      20'h04ca4: out <= 12'h000;
      20'h04ca5: out <= 12'h000;
      20'h04ca6: out <= 12'h000;
      20'h04ca7: out <= 12'h6af;
      20'h04ca8: out <= 12'h6af;
      20'h04ca9: out <= 12'h000;
      20'h04caa: out <= 12'h000;
      20'h04cab: out <= 12'h000;
      20'h04cac: out <= 12'h603;
      20'h04cad: out <= 12'h603;
      20'h04cae: out <= 12'h603;
      20'h04caf: out <= 12'h603;
      20'h04cb0: out <= 12'h222;
      20'h04cb1: out <= 12'h6af;
      20'h04cb2: out <= 12'h6af;
      20'h04cb3: out <= 12'h6af;
      20'h04cb4: out <= 12'h16d;
      20'h04cb5: out <= 12'h6af;
      20'h04cb6: out <= 12'h6af;
      20'h04cb7: out <= 12'h6af;
      20'h04cb8: out <= 12'h6af;
      20'h04cb9: out <= 12'h6af;
      20'h04cba: out <= 12'h6af;
      20'h04cbb: out <= 12'h6af;
      20'h04cbc: out <= 12'h6af;
      20'h04cbd: out <= 12'h6af;
      20'h04cbe: out <= 12'h6af;
      20'h04cbf: out <= 12'h6af;
      20'h04cc0: out <= 12'h603;
      20'h04cc1: out <= 12'h603;
      20'h04cc2: out <= 12'h603;
      20'h04cc3: out <= 12'h603;
      20'h04cc4: out <= 12'h000;
      20'h04cc5: out <= 12'h000;
      20'h04cc6: out <= 12'h16d;
      20'h04cc7: out <= 12'h6af;
      20'h04cc8: out <= 12'hfff;
      20'h04cc9: out <= 12'h6af;
      20'h04cca: out <= 12'h16d;
      20'h04ccb: out <= 12'h000;
      20'h04ccc: out <= 12'h603;
      20'h04ccd: out <= 12'h603;
      20'h04cce: out <= 12'h603;
      20'h04ccf: out <= 12'h603;
      20'h04cd0: out <= 12'h222;
      20'h04cd1: out <= 12'h222;
      20'h04cd2: out <= 12'h222;
      20'h04cd3: out <= 12'h660;
      20'h04cd4: out <= 12'h660;
      20'h04cd5: out <= 12'hbb0;
      20'h04cd6: out <= 12'hbb0;
      20'h04cd7: out <= 12'hbb0;
      20'h04cd8: out <= 12'hee9;
      20'h04cd9: out <= 12'hee9;
      20'h04cda: out <= 12'hee9;
      20'h04cdb: out <= 12'hee9;
      20'h04cdc: out <= 12'hee9;
      20'h04cdd: out <= 12'hbb0;
      20'h04cde: out <= 12'hbb0;
      20'h04cdf: out <= 12'h660;
      20'h04ce0: out <= 12'h603;
      20'h04ce1: out <= 12'h603;
      20'h04ce2: out <= 12'h603;
      20'h04ce3: out <= 12'h603;
      20'h04ce4: out <= 12'h000;
      20'h04ce5: out <= 12'h660;
      20'h04ce6: out <= 12'hbb0;
      20'h04ce7: out <= 12'hee9;
      20'h04ce8: out <= 12'hee9;
      20'h04ce9: out <= 12'hee9;
      20'h04cea: out <= 12'hbb0;
      20'h04ceb: out <= 12'h660;
      20'h04cec: out <= 12'h603;
      20'h04ced: out <= 12'h603;
      20'h04cee: out <= 12'h603;
      20'h04cef: out <= 12'h603;
      20'h04cf0: out <= 12'h222;
      20'h04cf1: out <= 12'h222;
      20'h04cf2: out <= 12'h222;
      20'h04cf3: out <= 12'h222;
      20'h04cf4: out <= 12'h222;
      20'h04cf5: out <= 12'h660;
      20'h04cf6: out <= 12'hbb0;
      20'h04cf7: out <= 12'hee9;
      20'h04cf8: out <= 12'hee9;
      20'h04cf9: out <= 12'hee9;
      20'h04cfa: out <= 12'hbb0;
      20'h04cfb: out <= 12'h660;
      20'h04cfc: out <= 12'h222;
      20'h04cfd: out <= 12'h222;
      20'h04cfe: out <= 12'h222;
      20'h04cff: out <= 12'h222;
      20'h04d00: out <= 12'h000;
      20'h04d01: out <= 12'h000;
      20'h04d02: out <= 12'h000;
      20'h04d03: out <= 12'h660;
      20'h04d04: out <= 12'hbb0;
      20'h04d05: out <= 12'hee9;
      20'h04d06: out <= 12'hee9;
      20'h04d07: out <= 12'hee9;
      20'h04d08: out <= 12'hee9;
      20'h04d09: out <= 12'hee9;
      20'h04d0a: out <= 12'hee9;
      20'h04d0b: out <= 12'hee9;
      20'h04d0c: out <= 12'hbb0;
      20'h04d0d: out <= 12'h660;
      20'h04d0e: out <= 12'h000;
      20'h04d0f: out <= 12'h000;
      20'h04d10: out <= 12'h603;
      20'h04d11: out <= 12'h603;
      20'h04d12: out <= 12'h603;
      20'h04d13: out <= 12'h603;
      20'h04d14: out <= 12'h000;
      20'h04d15: out <= 12'h666;
      20'h04d16: out <= 12'hfff;
      20'h04d17: out <= 12'h666;
      20'h04d18: out <= 12'h666;
      20'h04d19: out <= 12'hfff;
      20'h04d1a: out <= 12'h666;
      20'h04d1b: out <= 12'h666;
      20'h04d1c: out <= 12'h000;
      20'h04d1d: out <= 12'h666;
      20'h04d1e: out <= 12'h666;
      20'h04d1f: out <= 12'hfff;
      20'h04d20: out <= 12'h666;
      20'h04d21: out <= 12'h666;
      20'h04d22: out <= 12'hfff;
      20'h04d23: out <= 12'h666;
      20'h04d24: out <= 12'h000;
      20'h04d25: out <= 12'h000;
      20'h04d26: out <= 12'h000;
      20'h04d27: out <= 12'hb27;
      20'h04d28: out <= 12'hf87;
      20'h04d29: out <= 12'hee9;
      20'h04d2a: out <= 12'hee9;
      20'h04d2b: out <= 12'hf87;
      20'h04d2c: out <= 12'hf87;
      20'h04d2d: out <= 12'hf87;
      20'h04d2e: out <= 12'hb27;
      20'h04d2f: out <= 12'hb27;
      20'h04d30: out <= 12'hf87;
      20'h04d31: out <= 12'hee9;
      20'h04d32: out <= 12'h000;
      20'h04d33: out <= 12'h000;
      20'h04d34: out <= 12'h000;
      20'h04d35: out <= 12'h000;
      20'h04d36: out <= 12'h000;
      20'h04d37: out <= 12'hf87;
      20'h04d38: out <= 12'hf87;
      20'h04d39: out <= 12'hee9;
      20'h04d3a: out <= 12'hee9;
      20'h04d3b: out <= 12'hee9;
      20'h04d3c: out <= 12'hf87;
      20'h04d3d: out <= 12'hf87;
      20'h04d3e: out <= 12'hb27;
      20'h04d3f: out <= 12'hb27;
      20'h04d40: out <= 12'hb27;
      20'h04d41: out <= 12'hf87;
      20'h04d42: out <= 12'hf87;
      20'h04d43: out <= 12'h000;
      20'h04d44: out <= 12'h603;
      20'h04d45: out <= 12'h603;
      20'h04d46: out <= 12'h603;
      20'h04d47: out <= 12'h603;
      20'h04d48: out <= 12'h603;
      20'h04d49: out <= 12'h603;
      20'h04d4a: out <= 12'h603;
      20'h04d4b: out <= 12'h603;
      20'h04d4c: out <= 12'h603;
      20'h04d4d: out <= 12'h603;
      20'h04d4e: out <= 12'h603;
      20'h04d4f: out <= 12'h603;
      20'h04d50: out <= 12'h603;
      20'h04d51: out <= 12'h603;
      20'h04d52: out <= 12'h603;
      20'h04d53: out <= 12'h603;
      20'h04d54: out <= 12'h603;
      20'h04d55: out <= 12'h603;
      20'h04d56: out <= 12'h603;
      20'h04d57: out <= 12'h603;
      20'h04d58: out <= 12'h603;
      20'h04d59: out <= 12'h603;
      20'h04d5a: out <= 12'h603;
      20'h04d5b: out <= 12'h603;
      20'h04d5c: out <= 12'h603;
      20'h04d5d: out <= 12'h603;
      20'h04d5e: out <= 12'h603;
      20'h04d5f: out <= 12'h603;
      20'h04d60: out <= 12'h603;
      20'h04d61: out <= 12'h603;
      20'h04d62: out <= 12'h603;
      20'h04d63: out <= 12'h603;
      20'h04d64: out <= 12'h603;
      20'h04d65: out <= 12'h603;
      20'h04d66: out <= 12'h603;
      20'h04d67: out <= 12'h603;
      20'h04d68: out <= 12'hee9;
      20'h04d69: out <= 12'hf87;
      20'h04d6a: out <= 12'hf87;
      20'h04d6b: out <= 12'hf87;
      20'h04d6c: out <= 12'hf87;
      20'h04d6d: out <= 12'hf87;
      20'h04d6e: out <= 12'hf87;
      20'h04d6f: out <= 12'hb27;
      20'h04d70: out <= 12'h000;
      20'h04d71: out <= 12'h000;
      20'h04d72: out <= 12'h000;
      20'h04d73: out <= 12'h000;
      20'h04d74: out <= 12'h000;
      20'h04d75: out <= 12'h000;
      20'h04d76: out <= 12'h000;
      20'h04d77: out <= 12'h000;
      20'h04d78: out <= 12'h000;
      20'h04d79: out <= 12'h000;
      20'h04d7a: out <= 12'h000;
      20'h04d7b: out <= 12'h8d0;
      20'h04d7c: out <= 12'h8d0;
      20'h04d7d: out <= 12'h000;
      20'h04d7e: out <= 12'h000;
      20'h04d7f: out <= 12'h000;
      20'h04d80: out <= 12'h8d0;
      20'h04d81: out <= 12'h8d0;
      20'h04d82: out <= 12'h000;
      20'h04d83: out <= 12'h000;
      20'h04d84: out <= 12'h000;
      20'h04d85: out <= 12'h000;
      20'h04d86: out <= 12'h000;
      20'h04d87: out <= 12'h8d0;
      20'h04d88: out <= 12'h8d0;
      20'h04d89: out <= 12'h8d0;
      20'h04d8a: out <= 12'h8d0;
      20'h04d8b: out <= 12'h8d0;
      20'h04d8c: out <= 12'h000;
      20'h04d8d: out <= 12'h8d0;
      20'h04d8e: out <= 12'h8d0;
      20'h04d8f: out <= 12'h000;
      20'h04d90: out <= 12'h000;
      20'h04d91: out <= 12'h8d0;
      20'h04d92: out <= 12'h8d0;
      20'h04d93: out <= 12'h000;
      20'h04d94: out <= 12'h000;
      20'h04d95: out <= 12'h000;
      20'h04d96: out <= 12'h8d0;
      20'h04d97: out <= 12'h8d0;
      20'h04d98: out <= 12'h8d0;
      20'h04d99: out <= 12'h000;
      20'h04d9a: out <= 12'h000;
      20'h04d9b: out <= 12'h000;
      20'h04d9c: out <= 12'h000;
      20'h04d9d: out <= 12'h000;
      20'h04d9e: out <= 12'h000;
      20'h04d9f: out <= 12'h000;
      20'h04da0: out <= 12'h000;
      20'h04da1: out <= 12'h000;
      20'h04da2: out <= 12'h000;
      20'h04da3: out <= 12'h000;
      20'h04da4: out <= 12'h000;
      20'h04da5: out <= 12'h000;
      20'h04da6: out <= 12'h000;
      20'h04da7: out <= 12'h000;
      20'h04da8: out <= 12'h603;
      20'h04da9: out <= 12'h603;
      20'h04daa: out <= 12'h603;
      20'h04dab: out <= 12'h603;
      20'h04dac: out <= 12'h6af;
      20'h04dad: out <= 12'h6af;
      20'h04dae: out <= 12'h6af;
      20'h04daf: out <= 12'h6af;
      20'h04db0: out <= 12'h6af;
      20'h04db1: out <= 12'h6af;
      20'h04db2: out <= 12'h6af;
      20'h04db3: out <= 12'h6af;
      20'h04db4: out <= 12'h603;
      20'h04db5: out <= 12'h603;
      20'h04db6: out <= 12'h603;
      20'h04db7: out <= 12'h603;
      20'h04db8: out <= 12'h603;
      20'h04db9: out <= 12'h603;
      20'h04dba: out <= 12'h603;
      20'h04dbb: out <= 12'h603;
      20'h04dbc: out <= 12'h000;
      20'h04dbd: out <= 12'h000;
      20'h04dbe: out <= 12'h000;
      20'h04dbf: out <= 12'h6af;
      20'h04dc0: out <= 12'h6af;
      20'h04dc1: out <= 12'h000;
      20'h04dc2: out <= 12'h000;
      20'h04dc3: out <= 12'h000;
      20'h04dc4: out <= 12'h603;
      20'h04dc5: out <= 12'h603;
      20'h04dc6: out <= 12'h603;
      20'h04dc7: out <= 12'h603;
      20'h04dc8: out <= 12'h222;
      20'h04dc9: out <= 12'hfff;
      20'h04dca: out <= 12'hfff;
      20'h04dcb: out <= 12'hfff;
      20'h04dcc: out <= 12'h16d;
      20'h04dcd: out <= 12'hfff;
      20'h04dce: out <= 12'hfff;
      20'h04dcf: out <= 12'hfff;
      20'h04dd0: out <= 12'hfff;
      20'h04dd1: out <= 12'hfff;
      20'h04dd2: out <= 12'hfff;
      20'h04dd3: out <= 12'hfff;
      20'h04dd4: out <= 12'hfff;
      20'h04dd5: out <= 12'hfff;
      20'h04dd6: out <= 12'hfff;
      20'h04dd7: out <= 12'hfff;
      20'h04dd8: out <= 12'h603;
      20'h04dd9: out <= 12'h603;
      20'h04dda: out <= 12'h603;
      20'h04ddb: out <= 12'h603;
      20'h04ddc: out <= 12'h000;
      20'h04ddd: out <= 12'h000;
      20'h04dde: out <= 12'h16d;
      20'h04ddf: out <= 12'h6af;
      20'h04de0: out <= 12'hfff;
      20'h04de1: out <= 12'h6af;
      20'h04de2: out <= 12'h16d;
      20'h04de3: out <= 12'h000;
      20'h04de4: out <= 12'h603;
      20'h04de5: out <= 12'h603;
      20'h04de6: out <= 12'h603;
      20'h04de7: out <= 12'h603;
      20'h04de8: out <= 12'h660;
      20'h04de9: out <= 12'h660;
      20'h04dea: out <= 12'hbb0;
      20'h04deb: out <= 12'hbb0;
      20'h04dec: out <= 12'hbb0;
      20'h04ded: out <= 12'hee9;
      20'h04dee: out <= 12'hee9;
      20'h04def: out <= 12'hee9;
      20'h04df0: out <= 12'hee9;
      20'h04df1: out <= 12'hee9;
      20'h04df2: out <= 12'hee9;
      20'h04df3: out <= 12'hee9;
      20'h04df4: out <= 12'hee9;
      20'h04df5: out <= 12'hee9;
      20'h04df6: out <= 12'hee9;
      20'h04df7: out <= 12'hbb0;
      20'h04df8: out <= 12'h603;
      20'h04df9: out <= 12'h603;
      20'h04dfa: out <= 12'h603;
      20'h04dfb: out <= 12'h603;
      20'h04dfc: out <= 12'h000;
      20'h04dfd: out <= 12'h660;
      20'h04dfe: out <= 12'hbb0;
      20'h04dff: out <= 12'hee9;
      20'h04e00: out <= 12'hee9;
      20'h04e01: out <= 12'hee9;
      20'h04e02: out <= 12'hbb0;
      20'h04e03: out <= 12'h660;
      20'h04e04: out <= 12'h603;
      20'h04e05: out <= 12'h603;
      20'h04e06: out <= 12'h603;
      20'h04e07: out <= 12'h603;
      20'h04e08: out <= 12'h222;
      20'h04e09: out <= 12'h222;
      20'h04e0a: out <= 12'h222;
      20'h04e0b: out <= 12'h222;
      20'h04e0c: out <= 12'h222;
      20'h04e0d: out <= 12'h660;
      20'h04e0e: out <= 12'hbb0;
      20'h04e0f: out <= 12'hee9;
      20'h04e10: out <= 12'hee9;
      20'h04e11: out <= 12'hee9;
      20'h04e12: out <= 12'hbb0;
      20'h04e13: out <= 12'h660;
      20'h04e14: out <= 12'h222;
      20'h04e15: out <= 12'h222;
      20'h04e16: out <= 12'h222;
      20'h04e17: out <= 12'h222;
      20'h04e18: out <= 12'h000;
      20'h04e19: out <= 12'h660;
      20'h04e1a: out <= 12'hbb0;
      20'h04e1b: out <= 12'hee9;
      20'h04e1c: out <= 12'hee9;
      20'h04e1d: out <= 12'hee9;
      20'h04e1e: out <= 12'hee9;
      20'h04e1f: out <= 12'hee9;
      20'h04e20: out <= 12'hee9;
      20'h04e21: out <= 12'hee9;
      20'h04e22: out <= 12'hee9;
      20'h04e23: out <= 12'hee9;
      20'h04e24: out <= 12'hee9;
      20'h04e25: out <= 12'hee9;
      20'h04e26: out <= 12'hbb0;
      20'h04e27: out <= 12'h660;
      20'h04e28: out <= 12'h603;
      20'h04e29: out <= 12'h603;
      20'h04e2a: out <= 12'h603;
      20'h04e2b: out <= 12'h603;
      20'h04e2c: out <= 12'h000;
      20'h04e2d: out <= 12'h666;
      20'h04e2e: out <= 12'hfff;
      20'h04e2f: out <= 12'h666;
      20'h04e30: out <= 12'h666;
      20'h04e31: out <= 12'hfff;
      20'h04e32: out <= 12'h666;
      20'h04e33: out <= 12'h000;
      20'h04e34: out <= 12'h666;
      20'h04e35: out <= 12'h000;
      20'h04e36: out <= 12'h666;
      20'h04e37: out <= 12'hfff;
      20'h04e38: out <= 12'h666;
      20'h04e39: out <= 12'h666;
      20'h04e3a: out <= 12'hfff;
      20'h04e3b: out <= 12'h666;
      20'h04e3c: out <= 12'h000;
      20'h04e3d: out <= 12'h000;
      20'h04e3e: out <= 12'hb27;
      20'h04e3f: out <= 12'hf87;
      20'h04e40: out <= 12'hee9;
      20'h04e41: out <= 12'hf87;
      20'h04e42: out <= 12'hf87;
      20'h04e43: out <= 12'hb27;
      20'h04e44: out <= 12'hb27;
      20'h04e45: out <= 12'hb27;
      20'h04e46: out <= 12'hb27;
      20'h04e47: out <= 12'hb27;
      20'h04e48: out <= 12'hb27;
      20'h04e49: out <= 12'hb27;
      20'h04e4a: out <= 12'hee9;
      20'h04e4b: out <= 12'h000;
      20'h04e4c: out <= 12'h000;
      20'h04e4d: out <= 12'h000;
      20'h04e4e: out <= 12'h000;
      20'h04e4f: out <= 12'hb27;
      20'h04e50: out <= 12'hb27;
      20'h04e51: out <= 12'hb27;
      20'h04e52: out <= 12'hf87;
      20'h04e53: out <= 12'hf87;
      20'h04e54: out <= 12'hee9;
      20'h04e55: out <= 12'hb27;
      20'h04e56: out <= 12'hb27;
      20'h04e57: out <= 12'hb27;
      20'h04e58: out <= 12'hf87;
      20'h04e59: out <= 12'hf87;
      20'h04e5a: out <= 12'h000;
      20'h04e5b: out <= 12'h000;
      20'h04e5c: out <= 12'h603;
      20'h04e5d: out <= 12'h603;
      20'h04e5e: out <= 12'h603;
      20'h04e5f: out <= 12'h603;
      20'h04e60: out <= 12'h603;
      20'h04e61: out <= 12'h603;
      20'h04e62: out <= 12'h603;
      20'h04e63: out <= 12'h603;
      20'h04e64: out <= 12'h603;
      20'h04e65: out <= 12'h603;
      20'h04e66: out <= 12'h603;
      20'h04e67: out <= 12'h603;
      20'h04e68: out <= 12'h603;
      20'h04e69: out <= 12'h603;
      20'h04e6a: out <= 12'h603;
      20'h04e6b: out <= 12'h603;
      20'h04e6c: out <= 12'h603;
      20'h04e6d: out <= 12'h603;
      20'h04e6e: out <= 12'h603;
      20'h04e6f: out <= 12'h603;
      20'h04e70: out <= 12'h603;
      20'h04e71: out <= 12'h603;
      20'h04e72: out <= 12'h603;
      20'h04e73: out <= 12'h603;
      20'h04e74: out <= 12'h603;
      20'h04e75: out <= 12'h603;
      20'h04e76: out <= 12'h603;
      20'h04e77: out <= 12'h603;
      20'h04e78: out <= 12'h603;
      20'h04e79: out <= 12'h603;
      20'h04e7a: out <= 12'h603;
      20'h04e7b: out <= 12'h603;
      20'h04e7c: out <= 12'h603;
      20'h04e7d: out <= 12'h603;
      20'h04e7e: out <= 12'h603;
      20'h04e7f: out <= 12'h603;
      20'h04e80: out <= 12'hb27;
      20'h04e81: out <= 12'hb27;
      20'h04e82: out <= 12'hb27;
      20'h04e83: out <= 12'hb27;
      20'h04e84: out <= 12'hb27;
      20'h04e85: out <= 12'hb27;
      20'h04e86: out <= 12'hb27;
      20'h04e87: out <= 12'hb27;
      20'h04e88: out <= 12'h000;
      20'h04e89: out <= 12'h000;
      20'h04e8a: out <= 12'h000;
      20'h04e8b: out <= 12'h000;
      20'h04e8c: out <= 12'h000;
      20'h04e8d: out <= 12'h000;
      20'h04e8e: out <= 12'h000;
      20'h04e8f: out <= 12'h000;
      20'h04e90: out <= 12'h000;
      20'h04e91: out <= 12'h000;
      20'h04e92: out <= 12'h000;
      20'h04e93: out <= 12'h000;
      20'h04e94: out <= 12'h000;
      20'h04e95: out <= 12'h000;
      20'h04e96: out <= 12'h000;
      20'h04e97: out <= 12'h000;
      20'h04e98: out <= 12'h000;
      20'h04e99: out <= 12'h000;
      20'h04e9a: out <= 12'h000;
      20'h04e9b: out <= 12'h000;
      20'h04e9c: out <= 12'h000;
      20'h04e9d: out <= 12'h000;
      20'h04e9e: out <= 12'h000;
      20'h04e9f: out <= 12'h000;
      20'h04ea0: out <= 12'h000;
      20'h04ea1: out <= 12'h000;
      20'h04ea2: out <= 12'h000;
      20'h04ea3: out <= 12'h000;
      20'h04ea4: out <= 12'h000;
      20'h04ea5: out <= 12'h000;
      20'h04ea6: out <= 12'h000;
      20'h04ea7: out <= 12'h000;
      20'h04ea8: out <= 12'h000;
      20'h04ea9: out <= 12'h000;
      20'h04eaa: out <= 12'h000;
      20'h04eab: out <= 12'h000;
      20'h04eac: out <= 12'h000;
      20'h04ead: out <= 12'h000;
      20'h04eae: out <= 12'h000;
      20'h04eaf: out <= 12'h000;
      20'h04eb0: out <= 12'h000;
      20'h04eb1: out <= 12'h000;
      20'h04eb2: out <= 12'h000;
      20'h04eb3: out <= 12'h000;
      20'h04eb4: out <= 12'h000;
      20'h04eb5: out <= 12'h000;
      20'h04eb6: out <= 12'h000;
      20'h04eb7: out <= 12'h000;
      20'h04eb8: out <= 12'h000;
      20'h04eb9: out <= 12'h000;
      20'h04eba: out <= 12'h000;
      20'h04ebb: out <= 12'h000;
      20'h04ebc: out <= 12'h000;
      20'h04ebd: out <= 12'h000;
      20'h04ebe: out <= 12'h000;
      20'h04ebf: out <= 12'h000;
      20'h04ec0: out <= 12'h603;
      20'h04ec1: out <= 12'h603;
      20'h04ec2: out <= 12'h603;
      20'h04ec3: out <= 12'h603;
      20'h04ec4: out <= 12'h6af;
      20'h04ec5: out <= 12'h6af;
      20'h04ec6: out <= 12'h6af;
      20'h04ec7: out <= 12'h6af;
      20'h04ec8: out <= 12'h6af;
      20'h04ec9: out <= 12'h6af;
      20'h04eca: out <= 12'h6af;
      20'h04ecb: out <= 12'h6af;
      20'h04ecc: out <= 12'h603;
      20'h04ecd: out <= 12'h603;
      20'h04ece: out <= 12'h603;
      20'h04ecf: out <= 12'h603;
      20'h04ed0: out <= 12'h603;
      20'h04ed1: out <= 12'h603;
      20'h04ed2: out <= 12'h603;
      20'h04ed3: out <= 12'h603;
      20'h04ed4: out <= 12'h000;
      20'h04ed5: out <= 12'h000;
      20'h04ed6: out <= 12'h000;
      20'h04ed7: out <= 12'h6af;
      20'h04ed8: out <= 12'h6af;
      20'h04ed9: out <= 12'h000;
      20'h04eda: out <= 12'h000;
      20'h04edb: out <= 12'h000;
      20'h04edc: out <= 12'h603;
      20'h04edd: out <= 12'h603;
      20'h04ede: out <= 12'h603;
      20'h04edf: out <= 12'h603;
      20'h04ee0: out <= 12'h222;
      20'h04ee1: out <= 12'h6af;
      20'h04ee2: out <= 12'h6af;
      20'h04ee3: out <= 12'h6af;
      20'h04ee4: out <= 12'h16d;
      20'h04ee5: out <= 12'h6af;
      20'h04ee6: out <= 12'h6af;
      20'h04ee7: out <= 12'h6af;
      20'h04ee8: out <= 12'h6af;
      20'h04ee9: out <= 12'h6af;
      20'h04eea: out <= 12'h6af;
      20'h04eeb: out <= 12'h6af;
      20'h04eec: out <= 12'h6af;
      20'h04eed: out <= 12'h6af;
      20'h04eee: out <= 12'h6af;
      20'h04eef: out <= 12'h6af;
      20'h04ef0: out <= 12'h603;
      20'h04ef1: out <= 12'h603;
      20'h04ef2: out <= 12'h603;
      20'h04ef3: out <= 12'h603;
      20'h04ef4: out <= 12'h000;
      20'h04ef5: out <= 12'h000;
      20'h04ef6: out <= 12'h16d;
      20'h04ef7: out <= 12'h6af;
      20'h04ef8: out <= 12'hfff;
      20'h04ef9: out <= 12'h6af;
      20'h04efa: out <= 12'h16d;
      20'h04efb: out <= 12'h000;
      20'h04efc: out <= 12'h603;
      20'h04efd: out <= 12'h603;
      20'h04efe: out <= 12'h603;
      20'h04eff: out <= 12'h603;
      20'h04f00: out <= 12'h222;
      20'h04f01: out <= 12'h222;
      20'h04f02: out <= 12'h222;
      20'h04f03: out <= 12'h660;
      20'h04f04: out <= 12'h660;
      20'h04f05: out <= 12'hbb0;
      20'h04f06: out <= 12'hbb0;
      20'h04f07: out <= 12'hbb0;
      20'h04f08: out <= 12'hee9;
      20'h04f09: out <= 12'hee9;
      20'h04f0a: out <= 12'hee9;
      20'h04f0b: out <= 12'hee9;
      20'h04f0c: out <= 12'hee9;
      20'h04f0d: out <= 12'hbb0;
      20'h04f0e: out <= 12'hbb0;
      20'h04f0f: out <= 12'h660;
      20'h04f10: out <= 12'h603;
      20'h04f11: out <= 12'h603;
      20'h04f12: out <= 12'h603;
      20'h04f13: out <= 12'h603;
      20'h04f14: out <= 12'h000;
      20'h04f15: out <= 12'h000;
      20'h04f16: out <= 12'h660;
      20'h04f17: out <= 12'hbb0;
      20'h04f18: out <= 12'hee9;
      20'h04f19: out <= 12'hbb0;
      20'h04f1a: out <= 12'h660;
      20'h04f1b: out <= 12'h000;
      20'h04f1c: out <= 12'h603;
      20'h04f1d: out <= 12'h603;
      20'h04f1e: out <= 12'h603;
      20'h04f1f: out <= 12'h603;
      20'h04f20: out <= 12'h222;
      20'h04f21: out <= 12'h222;
      20'h04f22: out <= 12'h222;
      20'h04f23: out <= 12'h222;
      20'h04f24: out <= 12'h222;
      20'h04f25: out <= 12'h660;
      20'h04f26: out <= 12'hbb0;
      20'h04f27: out <= 12'hee9;
      20'h04f28: out <= 12'hee9;
      20'h04f29: out <= 12'hee9;
      20'h04f2a: out <= 12'hbb0;
      20'h04f2b: out <= 12'h660;
      20'h04f2c: out <= 12'h222;
      20'h04f2d: out <= 12'h222;
      20'h04f2e: out <= 12'h222;
      20'h04f2f: out <= 12'h222;
      20'h04f30: out <= 12'h000;
      20'h04f31: out <= 12'h000;
      20'h04f32: out <= 12'h000;
      20'h04f33: out <= 12'h660;
      20'h04f34: out <= 12'hbb0;
      20'h04f35: out <= 12'hee9;
      20'h04f36: out <= 12'hee9;
      20'h04f37: out <= 12'hee9;
      20'h04f38: out <= 12'hee9;
      20'h04f39: out <= 12'hee9;
      20'h04f3a: out <= 12'hee9;
      20'h04f3b: out <= 12'hee9;
      20'h04f3c: out <= 12'hbb0;
      20'h04f3d: out <= 12'h660;
      20'h04f3e: out <= 12'h000;
      20'h04f3f: out <= 12'h000;
      20'h04f40: out <= 12'h603;
      20'h04f41: out <= 12'h603;
      20'h04f42: out <= 12'h603;
      20'h04f43: out <= 12'h603;
      20'h04f44: out <= 12'h000;
      20'h04f45: out <= 12'h666;
      20'h04f46: out <= 12'hfff;
      20'h04f47: out <= 12'h666;
      20'h04f48: out <= 12'h666;
      20'h04f49: out <= 12'hfff;
      20'h04f4a: out <= 12'h000;
      20'h04f4b: out <= 12'h666;
      20'h04f4c: out <= 12'h666;
      20'h04f4d: out <= 12'h666;
      20'h04f4e: out <= 12'h000;
      20'h04f4f: out <= 12'hfff;
      20'h04f50: out <= 12'h666;
      20'h04f51: out <= 12'h666;
      20'h04f52: out <= 12'hfff;
      20'h04f53: out <= 12'h666;
      20'h04f54: out <= 12'h000;
      20'h04f55: out <= 12'h000;
      20'h04f56: out <= 12'h000;
      20'h04f57: out <= 12'hb27;
      20'h04f58: out <= 12'hf87;
      20'h04f59: out <= 12'hee9;
      20'h04f5a: out <= 12'hee9;
      20'h04f5b: out <= 12'hf87;
      20'h04f5c: out <= 12'hf87;
      20'h04f5d: out <= 12'hf87;
      20'h04f5e: out <= 12'hb27;
      20'h04f5f: out <= 12'hb27;
      20'h04f60: out <= 12'hf87;
      20'h04f61: out <= 12'hee9;
      20'h04f62: out <= 12'h000;
      20'h04f63: out <= 12'h000;
      20'h04f64: out <= 12'h000;
      20'h04f65: out <= 12'h000;
      20'h04f66: out <= 12'h000;
      20'h04f67: out <= 12'h000;
      20'h04f68: out <= 12'hb27;
      20'h04f69: out <= 12'hf87;
      20'h04f6a: out <= 12'hb27;
      20'h04f6b: out <= 12'hb27;
      20'h04f6c: out <= 12'hb27;
      20'h04f6d: out <= 12'hee9;
      20'h04f6e: out <= 12'hf87;
      20'h04f6f: out <= 12'hf87;
      20'h04f70: out <= 12'hee9;
      20'h04f71: out <= 12'hf87;
      20'h04f72: out <= 12'h000;
      20'h04f73: out <= 12'h000;
      20'h04f74: out <= 12'h603;
      20'h04f75: out <= 12'h603;
      20'h04f76: out <= 12'h603;
      20'h04f77: out <= 12'h603;
      20'h04f78: out <= 12'h603;
      20'h04f79: out <= 12'h603;
      20'h04f7a: out <= 12'h603;
      20'h04f7b: out <= 12'h603;
      20'h04f7c: out <= 12'h603;
      20'h04f7d: out <= 12'h603;
      20'h04f7e: out <= 12'h603;
      20'h04f7f: out <= 12'h603;
      20'h04f80: out <= 12'h603;
      20'h04f81: out <= 12'h603;
      20'h04f82: out <= 12'h603;
      20'h04f83: out <= 12'h603;
      20'h04f84: out <= 12'h603;
      20'h04f85: out <= 12'h603;
      20'h04f86: out <= 12'h603;
      20'h04f87: out <= 12'h603;
      20'h04f88: out <= 12'h603;
      20'h04f89: out <= 12'h603;
      20'h04f8a: out <= 12'h603;
      20'h04f8b: out <= 12'h603;
      20'h04f8c: out <= 12'h603;
      20'h04f8d: out <= 12'h603;
      20'h04f8e: out <= 12'h603;
      20'h04f8f: out <= 12'h603;
      20'h04f90: out <= 12'h603;
      20'h04f91: out <= 12'h603;
      20'h04f92: out <= 12'h603;
      20'h04f93: out <= 12'h603;
      20'h04f94: out <= 12'h603;
      20'h04f95: out <= 12'h603;
      20'h04f96: out <= 12'h603;
      20'h04f97: out <= 12'h603;
      20'h04f98: out <= 12'hee9;
      20'h04f99: out <= 12'hee9;
      20'h04f9a: out <= 12'hee9;
      20'h04f9b: out <= 12'hee9;
      20'h04f9c: out <= 12'hee9;
      20'h04f9d: out <= 12'hee9;
      20'h04f9e: out <= 12'hee9;
      20'h04f9f: out <= 12'hb27;
      20'h04fa0: out <= 12'h000;
      20'h04fa1: out <= 12'h000;
      20'h04fa2: out <= 12'h000;
      20'h04fa3: out <= 12'h000;
      20'h04fa4: out <= 12'h000;
      20'h04fa5: out <= 12'h000;
      20'h04fa6: out <= 12'h000;
      20'h04fa7: out <= 12'h000;
      20'h04fa8: out <= 12'h000;
      20'h04fa9: out <= 12'h000;
      20'h04faa: out <= 12'h000;
      20'h04fab: out <= 12'h000;
      20'h04fac: out <= 12'h000;
      20'h04fad: out <= 12'h000;
      20'h04fae: out <= 12'h000;
      20'h04faf: out <= 12'h6af;
      20'h04fb0: out <= 12'hfff;
      20'h04fb1: out <= 12'h6af;
      20'h04fb2: out <= 12'h000;
      20'h04fb3: out <= 12'h000;
      20'h04fb4: out <= 12'h000;
      20'h04fb5: out <= 12'h000;
      20'h04fb6: out <= 12'h000;
      20'h04fb7: out <= 12'h000;
      20'h04fb8: out <= 12'h000;
      20'h04fb9: out <= 12'h000;
      20'h04fba: out <= 12'h000;
      20'h04fbb: out <= 12'h000;
      20'h04fbc: out <= 12'h000;
      20'h04fbd: out <= 12'h000;
      20'h04fbe: out <= 12'h000;
      20'h04fbf: out <= 12'h000;
      20'h04fc0: out <= 12'h000;
      20'h04fc1: out <= 12'h000;
      20'h04fc2: out <= 12'h000;
      20'h04fc3: out <= 12'h000;
      20'h04fc4: out <= 12'h000;
      20'h04fc5: out <= 12'h000;
      20'h04fc6: out <= 12'h000;
      20'h04fc7: out <= 12'h000;
      20'h04fc8: out <= 12'h000;
      20'h04fc9: out <= 12'h000;
      20'h04fca: out <= 12'h000;
      20'h04fcb: out <= 12'h000;
      20'h04fcc: out <= 12'h000;
      20'h04fcd: out <= 12'h000;
      20'h04fce: out <= 12'h000;
      20'h04fcf: out <= 12'h000;
      20'h04fd0: out <= 12'h000;
      20'h04fd1: out <= 12'h000;
      20'h04fd2: out <= 12'h000;
      20'h04fd3: out <= 12'h000;
      20'h04fd4: out <= 12'h000;
      20'h04fd5: out <= 12'h000;
      20'h04fd6: out <= 12'h000;
      20'h04fd7: out <= 12'h000;
      20'h04fd8: out <= 12'h603;
      20'h04fd9: out <= 12'h603;
      20'h04fda: out <= 12'h603;
      20'h04fdb: out <= 12'h603;
      20'h04fdc: out <= 12'h222;
      20'h04fdd: out <= 12'h222;
      20'h04fde: out <= 12'h222;
      20'h04fdf: out <= 12'h222;
      20'h04fe0: out <= 12'h222;
      20'h04fe1: out <= 12'h222;
      20'h04fe2: out <= 12'h222;
      20'h04fe3: out <= 12'h222;
      20'h04fe4: out <= 12'h603;
      20'h04fe5: out <= 12'h603;
      20'h04fe6: out <= 12'h603;
      20'h04fe7: out <= 12'h603;
      20'h04fe8: out <= 12'h603;
      20'h04fe9: out <= 12'h603;
      20'h04fea: out <= 12'h603;
      20'h04feb: out <= 12'h603;
      20'h04fec: out <= 12'h000;
      20'h04fed: out <= 12'h000;
      20'h04fee: out <= 12'h000;
      20'h04fef: out <= 12'h6af;
      20'h04ff0: out <= 12'h6af;
      20'h04ff1: out <= 12'h000;
      20'h04ff2: out <= 12'h000;
      20'h04ff3: out <= 12'h000;
      20'h04ff4: out <= 12'h603;
      20'h04ff5: out <= 12'h603;
      20'h04ff6: out <= 12'h603;
      20'h04ff7: out <= 12'h603;
      20'h04ff8: out <= 12'h222;
      20'h04ff9: out <= 12'h16d;
      20'h04ffa: out <= 12'h16d;
      20'h04ffb: out <= 12'h16d;
      20'h04ffc: out <= 12'h222;
      20'h04ffd: out <= 12'h16d;
      20'h04ffe: out <= 12'h16d;
      20'h04fff: out <= 12'h16d;
      20'h05000: out <= 12'h16d;
      20'h05001: out <= 12'h16d;
      20'h05002: out <= 12'h16d;
      20'h05003: out <= 12'h16d;
      20'h05004: out <= 12'h16d;
      20'h05005: out <= 12'h16d;
      20'h05006: out <= 12'h16d;
      20'h05007: out <= 12'h222;
      20'h05008: out <= 12'h603;
      20'h05009: out <= 12'h603;
      20'h0500a: out <= 12'h603;
      20'h0500b: out <= 12'h603;
      20'h0500c: out <= 12'h000;
      20'h0500d: out <= 12'h000;
      20'h0500e: out <= 12'h16d;
      20'h0500f: out <= 12'h6af;
      20'h05010: out <= 12'hfff;
      20'h05011: out <= 12'h6af;
      20'h05012: out <= 12'h16d;
      20'h05013: out <= 12'h000;
      20'h05014: out <= 12'h603;
      20'h05015: out <= 12'h603;
      20'h05016: out <= 12'h603;
      20'h05017: out <= 12'h603;
      20'h05018: out <= 12'h222;
      20'h05019: out <= 12'h222;
      20'h0501a: out <= 12'h222;
      20'h0501b: out <= 12'h222;
      20'h0501c: out <= 12'h222;
      20'h0501d: out <= 12'h222;
      20'h0501e: out <= 12'h660;
      20'h0501f: out <= 12'h660;
      20'h05020: out <= 12'hbb0;
      20'h05021: out <= 12'hbb0;
      20'h05022: out <= 12'hbb0;
      20'h05023: out <= 12'hbb0;
      20'h05024: out <= 12'hbb0;
      20'h05025: out <= 12'h660;
      20'h05026: out <= 12'h660;
      20'h05027: out <= 12'h222;
      20'h05028: out <= 12'h603;
      20'h05029: out <= 12'h603;
      20'h0502a: out <= 12'h603;
      20'h0502b: out <= 12'h603;
      20'h0502c: out <= 12'h000;
      20'h0502d: out <= 12'h000;
      20'h0502e: out <= 12'h660;
      20'h0502f: out <= 12'hbb0;
      20'h05030: out <= 12'hee9;
      20'h05031: out <= 12'hbb0;
      20'h05032: out <= 12'h660;
      20'h05033: out <= 12'h000;
      20'h05034: out <= 12'h603;
      20'h05035: out <= 12'h603;
      20'h05036: out <= 12'h603;
      20'h05037: out <= 12'h603;
      20'h05038: out <= 12'h222;
      20'h05039: out <= 12'h222;
      20'h0503a: out <= 12'h222;
      20'h0503b: out <= 12'h222;
      20'h0503c: out <= 12'h222;
      20'h0503d: out <= 12'h222;
      20'h0503e: out <= 12'hee9;
      20'h0503f: out <= 12'hbb0;
      20'h05040: out <= 12'hbb0;
      20'h05041: out <= 12'hbb0;
      20'h05042: out <= 12'hee9;
      20'h05043: out <= 12'h222;
      20'h05044: out <= 12'h222;
      20'h05045: out <= 12'h222;
      20'h05046: out <= 12'h222;
      20'h05047: out <= 12'h222;
      20'h05048: out <= 12'h000;
      20'h05049: out <= 12'h000;
      20'h0504a: out <= 12'h000;
      20'h0504b: out <= 12'h000;
      20'h0504c: out <= 12'h660;
      20'h0504d: out <= 12'hbb0;
      20'h0504e: out <= 12'hee9;
      20'h0504f: out <= 12'hee9;
      20'h05050: out <= 12'hee9;
      20'h05051: out <= 12'hee9;
      20'h05052: out <= 12'hee9;
      20'h05053: out <= 12'hbb0;
      20'h05054: out <= 12'h660;
      20'h05055: out <= 12'h000;
      20'h05056: out <= 12'h000;
      20'h05057: out <= 12'h000;
      20'h05058: out <= 12'h603;
      20'h05059: out <= 12'h603;
      20'h0505a: out <= 12'h603;
      20'h0505b: out <= 12'h603;
      20'h0505c: out <= 12'h000;
      20'h0505d: out <= 12'h666;
      20'h0505e: out <= 12'hfff;
      20'h0505f: out <= 12'h666;
      20'h05060: out <= 12'h666;
      20'h05061: out <= 12'h000;
      20'h05062: out <= 12'hfff;
      20'h05063: out <= 12'hfff;
      20'h05064: out <= 12'hfff;
      20'h05065: out <= 12'hfff;
      20'h05066: out <= 12'hfff;
      20'h05067: out <= 12'h000;
      20'h05068: out <= 12'h666;
      20'h05069: out <= 12'h666;
      20'h0506a: out <= 12'hfff;
      20'h0506b: out <= 12'h666;
      20'h0506c: out <= 12'h000;
      20'h0506d: out <= 12'h000;
      20'h0506e: out <= 12'h000;
      20'h0506f: out <= 12'hb27;
      20'h05070: out <= 12'hf87;
      20'h05071: out <= 12'hee9;
      20'h05072: out <= 12'hee9;
      20'h05073: out <= 12'hf87;
      20'h05074: out <= 12'hf87;
      20'h05075: out <= 12'hf87;
      20'h05076: out <= 12'hb27;
      20'h05077: out <= 12'hb27;
      20'h05078: out <= 12'hf87;
      20'h05079: out <= 12'hee9;
      20'h0507a: out <= 12'h000;
      20'h0507b: out <= 12'h000;
      20'h0507c: out <= 12'h000;
      20'h0507d: out <= 12'h000;
      20'h0507e: out <= 12'h000;
      20'h0507f: out <= 12'h000;
      20'h05080: out <= 12'hb27;
      20'h05081: out <= 12'hf87;
      20'h05082: out <= 12'hee9;
      20'h05083: out <= 12'hee9;
      20'h05084: out <= 12'hf87;
      20'h05085: out <= 12'hb27;
      20'h05086: out <= 12'hb27;
      20'h05087: out <= 12'hb27;
      20'h05088: out <= 12'hb27;
      20'h05089: out <= 12'hee9;
      20'h0508a: out <= 12'hee9;
      20'h0508b: out <= 12'h000;
      20'h0508c: out <= 12'h603;
      20'h0508d: out <= 12'h603;
      20'h0508e: out <= 12'h603;
      20'h0508f: out <= 12'h603;
      20'h05090: out <= 12'h603;
      20'h05091: out <= 12'h603;
      20'h05092: out <= 12'h603;
      20'h05093: out <= 12'h603;
      20'h05094: out <= 12'h603;
      20'h05095: out <= 12'h603;
      20'h05096: out <= 12'h603;
      20'h05097: out <= 12'h603;
      20'h05098: out <= 12'h603;
      20'h05099: out <= 12'h603;
      20'h0509a: out <= 12'h603;
      20'h0509b: out <= 12'h603;
      20'h0509c: out <= 12'h603;
      20'h0509d: out <= 12'h603;
      20'h0509e: out <= 12'h603;
      20'h0509f: out <= 12'h603;
      20'h050a0: out <= 12'h603;
      20'h050a1: out <= 12'h603;
      20'h050a2: out <= 12'h603;
      20'h050a3: out <= 12'h603;
      20'h050a4: out <= 12'h603;
      20'h050a5: out <= 12'h603;
      20'h050a6: out <= 12'h603;
      20'h050a7: out <= 12'h603;
      20'h050a8: out <= 12'h603;
      20'h050a9: out <= 12'h603;
      20'h050aa: out <= 12'h603;
      20'h050ab: out <= 12'h603;
      20'h050ac: out <= 12'h603;
      20'h050ad: out <= 12'h603;
      20'h050ae: out <= 12'h603;
      20'h050af: out <= 12'h603;
      20'h050b0: out <= 12'hee9;
      20'h050b1: out <= 12'hf87;
      20'h050b2: out <= 12'hf87;
      20'h050b3: out <= 12'hf87;
      20'h050b4: out <= 12'hf87;
      20'h050b5: out <= 12'hf87;
      20'h050b6: out <= 12'hf87;
      20'h050b7: out <= 12'hb27;
      20'h050b8: out <= 12'h000;
      20'h050b9: out <= 12'h000;
      20'h050ba: out <= 12'h000;
      20'h050bb: out <= 12'h000;
      20'h050bc: out <= 12'h000;
      20'h050bd: out <= 12'h000;
      20'h050be: out <= 12'h000;
      20'h050bf: out <= 12'h000;
      20'h050c0: out <= 12'h000;
      20'h050c1: out <= 12'h000;
      20'h050c2: out <= 12'h000;
      20'h050c3: out <= 12'h000;
      20'h050c4: out <= 12'h000;
      20'h050c5: out <= 12'h000;
      20'h050c6: out <= 12'h000;
      20'h050c7: out <= 12'h16d;
      20'h050c8: out <= 12'hfff;
      20'h050c9: out <= 12'h16d;
      20'h050ca: out <= 12'h000;
      20'h050cb: out <= 12'h000;
      20'h050cc: out <= 12'h000;
      20'h050cd: out <= 12'h000;
      20'h050ce: out <= 12'h000;
      20'h050cf: out <= 12'h000;
      20'h050d0: out <= 12'h000;
      20'h050d1: out <= 12'h000;
      20'h050d2: out <= 12'h000;
      20'h050d3: out <= 12'h000;
      20'h050d4: out <= 12'h000;
      20'h050d5: out <= 12'h000;
      20'h050d6: out <= 12'h000;
      20'h050d7: out <= 12'h000;
      20'h050d8: out <= 12'h000;
      20'h050d9: out <= 12'h000;
      20'h050da: out <= 12'h000;
      20'h050db: out <= 12'h000;
      20'h050dc: out <= 12'h000;
      20'h050dd: out <= 12'h000;
      20'h050de: out <= 12'h000;
      20'h050df: out <= 12'h000;
      20'h050e0: out <= 12'h000;
      20'h050e1: out <= 12'h000;
      20'h050e2: out <= 12'h000;
      20'h050e3: out <= 12'h000;
      20'h050e4: out <= 12'h000;
      20'h050e5: out <= 12'h000;
      20'h050e6: out <= 12'h000;
      20'h050e7: out <= 12'h000;
      20'h050e8: out <= 12'h000;
      20'h050e9: out <= 12'h000;
      20'h050ea: out <= 12'h000;
      20'h050eb: out <= 12'h000;
      20'h050ec: out <= 12'h000;
      20'h050ed: out <= 12'h000;
      20'h050ee: out <= 12'h000;
      20'h050ef: out <= 12'h000;
      20'h050f0: out <= 12'h603;
      20'h050f1: out <= 12'h603;
      20'h050f2: out <= 12'h603;
      20'h050f3: out <= 12'h603;
      20'h050f4: out <= 12'h222;
      20'h050f5: out <= 12'h222;
      20'h050f6: out <= 12'h222;
      20'h050f7: out <= 12'h222;
      20'h050f8: out <= 12'h222;
      20'h050f9: out <= 12'h222;
      20'h050fa: out <= 12'h222;
      20'h050fb: out <= 12'h222;
      20'h050fc: out <= 12'h603;
      20'h050fd: out <= 12'h603;
      20'h050fe: out <= 12'h603;
      20'h050ff: out <= 12'h603;
      20'h05100: out <= 12'h603;
      20'h05101: out <= 12'h603;
      20'h05102: out <= 12'h603;
      20'h05103: out <= 12'h603;
      20'h05104: out <= 12'h000;
      20'h05105: out <= 12'h000;
      20'h05106: out <= 12'h000;
      20'h05107: out <= 12'h6af;
      20'h05108: out <= 12'h6af;
      20'h05109: out <= 12'h000;
      20'h0510a: out <= 12'h000;
      20'h0510b: out <= 12'h000;
      20'h0510c: out <= 12'h603;
      20'h0510d: out <= 12'h603;
      20'h0510e: out <= 12'h603;
      20'h0510f: out <= 12'h603;
      20'h05110: out <= 12'h222;
      20'h05111: out <= 12'h6af;
      20'h05112: out <= 12'h6af;
      20'h05113: out <= 12'h222;
      20'h05114: out <= 12'h222;
      20'h05115: out <= 12'h222;
      20'h05116: out <= 12'h222;
      20'h05117: out <= 12'h222;
      20'h05118: out <= 12'h222;
      20'h05119: out <= 12'h222;
      20'h0511a: out <= 12'h222;
      20'h0511b: out <= 12'h222;
      20'h0511c: out <= 12'h222;
      20'h0511d: out <= 12'h222;
      20'h0511e: out <= 12'h222;
      20'h0511f: out <= 12'h222;
      20'h05120: out <= 12'h603;
      20'h05121: out <= 12'h603;
      20'h05122: out <= 12'h603;
      20'h05123: out <= 12'h603;
      20'h05124: out <= 12'h000;
      20'h05125: out <= 12'h000;
      20'h05126: out <= 12'h16d;
      20'h05127: out <= 12'h6af;
      20'h05128: out <= 12'hfff;
      20'h05129: out <= 12'h6af;
      20'h0512a: out <= 12'h16d;
      20'h0512b: out <= 12'h000;
      20'h0512c: out <= 12'h603;
      20'h0512d: out <= 12'h603;
      20'h0512e: out <= 12'h603;
      20'h0512f: out <= 12'h603;
      20'h05130: out <= 12'h222;
      20'h05131: out <= 12'h222;
      20'h05132: out <= 12'h222;
      20'h05133: out <= 12'h222;
      20'h05134: out <= 12'h222;
      20'h05135: out <= 12'h222;
      20'h05136: out <= 12'h222;
      20'h05137: out <= 12'h222;
      20'h05138: out <= 12'h660;
      20'h05139: out <= 12'h660;
      20'h0513a: out <= 12'h660;
      20'h0513b: out <= 12'h660;
      20'h0513c: out <= 12'h660;
      20'h0513d: out <= 12'h222;
      20'h0513e: out <= 12'h222;
      20'h0513f: out <= 12'h222;
      20'h05140: out <= 12'h603;
      20'h05141: out <= 12'h603;
      20'h05142: out <= 12'h603;
      20'h05143: out <= 12'h603;
      20'h05144: out <= 12'h000;
      20'h05145: out <= 12'h000;
      20'h05146: out <= 12'h000;
      20'h05147: out <= 12'hbb0;
      20'h05148: out <= 12'hee9;
      20'h05149: out <= 12'hbb0;
      20'h0514a: out <= 12'h000;
      20'h0514b: out <= 12'h000;
      20'h0514c: out <= 12'h603;
      20'h0514d: out <= 12'h603;
      20'h0514e: out <= 12'h603;
      20'h0514f: out <= 12'h603;
      20'h05150: out <= 12'h222;
      20'h05151: out <= 12'h222;
      20'h05152: out <= 12'h222;
      20'h05153: out <= 12'h222;
      20'h05154: out <= 12'h222;
      20'h05155: out <= 12'hbb0;
      20'h05156: out <= 12'h222;
      20'h05157: out <= 12'h660;
      20'h05158: out <= 12'h660;
      20'h05159: out <= 12'h660;
      20'h0515a: out <= 12'h222;
      20'h0515b: out <= 12'hbb0;
      20'h0515c: out <= 12'h222;
      20'h0515d: out <= 12'h222;
      20'h0515e: out <= 12'h222;
      20'h0515f: out <= 12'h222;
      20'h05160: out <= 12'h000;
      20'h05161: out <= 12'h000;
      20'h05162: out <= 12'h000;
      20'h05163: out <= 12'h000;
      20'h05164: out <= 12'h000;
      20'h05165: out <= 12'h660;
      20'h05166: out <= 12'hbb0;
      20'h05167: out <= 12'hee9;
      20'h05168: out <= 12'hee9;
      20'h05169: out <= 12'hee9;
      20'h0516a: out <= 12'hbb0;
      20'h0516b: out <= 12'h660;
      20'h0516c: out <= 12'h000;
      20'h0516d: out <= 12'h000;
      20'h0516e: out <= 12'h000;
      20'h0516f: out <= 12'h000;
      20'h05170: out <= 12'h603;
      20'h05171: out <= 12'h603;
      20'h05172: out <= 12'h603;
      20'h05173: out <= 12'h603;
      20'h05174: out <= 12'h000;
      20'h05175: out <= 12'h666;
      20'h05176: out <= 12'hfff;
      20'h05177: out <= 12'hfff;
      20'h05178: out <= 12'h000;
      20'h05179: out <= 12'hfff;
      20'h0517a: out <= 12'hfff;
      20'h0517b: out <= 12'hfff;
      20'h0517c: out <= 12'hfff;
      20'h0517d: out <= 12'hfff;
      20'h0517e: out <= 12'hfff;
      20'h0517f: out <= 12'hfff;
      20'h05180: out <= 12'h000;
      20'h05181: out <= 12'hfff;
      20'h05182: out <= 12'hfff;
      20'h05183: out <= 12'h666;
      20'h05184: out <= 12'h000;
      20'h05185: out <= 12'h000;
      20'h05186: out <= 12'h000;
      20'h05187: out <= 12'hb27;
      20'h05188: out <= 12'hf87;
      20'h05189: out <= 12'hee9;
      20'h0518a: out <= 12'hee9;
      20'h0518b: out <= 12'hf87;
      20'h0518c: out <= 12'hf87;
      20'h0518d: out <= 12'hf87;
      20'h0518e: out <= 12'hb27;
      20'h0518f: out <= 12'hb27;
      20'h05190: out <= 12'hf87;
      20'h05191: out <= 12'hee9;
      20'h05192: out <= 12'h000;
      20'h05193: out <= 12'h000;
      20'h05194: out <= 12'h000;
      20'h05195: out <= 12'h000;
      20'h05196: out <= 12'h000;
      20'h05197: out <= 12'h000;
      20'h05198: out <= 12'hb27;
      20'h05199: out <= 12'hf87;
      20'h0519a: out <= 12'hf87;
      20'h0519b: out <= 12'hee9;
      20'h0519c: out <= 12'hee9;
      20'h0519d: out <= 12'hf87;
      20'h0519e: out <= 12'hb27;
      20'h0519f: out <= 12'hb27;
      20'h051a0: out <= 12'hf87;
      20'h051a1: out <= 12'hb27;
      20'h051a2: out <= 12'h000;
      20'h051a3: out <= 12'h000;
      20'h051a4: out <= 12'h603;
      20'h051a5: out <= 12'h603;
      20'h051a6: out <= 12'h603;
      20'h051a7: out <= 12'h603;
      20'h051a8: out <= 12'h603;
      20'h051a9: out <= 12'h603;
      20'h051aa: out <= 12'h603;
      20'h051ab: out <= 12'h603;
      20'h051ac: out <= 12'h603;
      20'h051ad: out <= 12'h603;
      20'h051ae: out <= 12'h603;
      20'h051af: out <= 12'h603;
      20'h051b0: out <= 12'h603;
      20'h051b1: out <= 12'h603;
      20'h051b2: out <= 12'h603;
      20'h051b3: out <= 12'h603;
      20'h051b4: out <= 12'h603;
      20'h051b5: out <= 12'h603;
      20'h051b6: out <= 12'h603;
      20'h051b7: out <= 12'h603;
      20'h051b8: out <= 12'h603;
      20'h051b9: out <= 12'h603;
      20'h051ba: out <= 12'h603;
      20'h051bb: out <= 12'h603;
      20'h051bc: out <= 12'h603;
      20'h051bd: out <= 12'h603;
      20'h051be: out <= 12'h603;
      20'h051bf: out <= 12'h603;
      20'h051c0: out <= 12'h603;
      20'h051c1: out <= 12'h603;
      20'h051c2: out <= 12'h603;
      20'h051c3: out <= 12'h603;
      20'h051c4: out <= 12'h603;
      20'h051c5: out <= 12'h603;
      20'h051c6: out <= 12'h603;
      20'h051c7: out <= 12'h603;
      20'h051c8: out <= 12'hee9;
      20'h051c9: out <= 12'hf87;
      20'h051ca: out <= 12'hee9;
      20'h051cb: out <= 12'hee9;
      20'h051cc: out <= 12'hee9;
      20'h051cd: out <= 12'hb27;
      20'h051ce: out <= 12'hf87;
      20'h051cf: out <= 12'hb27;
      20'h051d0: out <= 12'h000;
      20'h051d1: out <= 12'h000;
      20'h051d2: out <= 12'h000;
      20'h051d3: out <= 12'h000;
      20'h051d4: out <= 12'h000;
      20'h051d5: out <= 12'h000;
      20'h051d6: out <= 12'h000;
      20'h051d7: out <= 12'h000;
      20'h051d8: out <= 12'h000;
      20'h051d9: out <= 12'h000;
      20'h051da: out <= 12'h000;
      20'h051db: out <= 12'h000;
      20'h051dc: out <= 12'h000;
      20'h051dd: out <= 12'h000;
      20'h051de: out <= 12'h000;
      20'h051df: out <= 12'h16d;
      20'h051e0: out <= 12'hfff;
      20'h051e1: out <= 12'h16d;
      20'h051e2: out <= 12'h000;
      20'h051e3: out <= 12'h000;
      20'h051e4: out <= 12'h000;
      20'h051e5: out <= 12'h000;
      20'h051e6: out <= 12'h000;
      20'h051e7: out <= 12'h000;
      20'h051e8: out <= 12'h000;
      20'h051e9: out <= 12'h000;
      20'h051ea: out <= 12'h000;
      20'h051eb: out <= 12'h000;
      20'h051ec: out <= 12'h000;
      20'h051ed: out <= 12'h000;
      20'h051ee: out <= 12'h000;
      20'h051ef: out <= 12'h000;
      20'h051f0: out <= 12'h000;
      20'h051f1: out <= 12'h000;
      20'h051f2: out <= 12'h000;
      20'h051f3: out <= 12'h000;
      20'h051f4: out <= 12'h000;
      20'h051f5: out <= 12'h000;
      20'h051f6: out <= 12'h000;
      20'h051f7: out <= 12'h000;
      20'h051f8: out <= 12'h000;
      20'h051f9: out <= 12'h000;
      20'h051fa: out <= 12'h000;
      20'h051fb: out <= 12'h000;
      20'h051fc: out <= 12'h000;
      20'h051fd: out <= 12'h000;
      20'h051fe: out <= 12'h000;
      20'h051ff: out <= 12'h000;
      20'h05200: out <= 12'h000;
      20'h05201: out <= 12'h000;
      20'h05202: out <= 12'h000;
      20'h05203: out <= 12'h000;
      20'h05204: out <= 12'h000;
      20'h05205: out <= 12'h000;
      20'h05206: out <= 12'h000;
      20'h05207: out <= 12'h000;
      20'h05208: out <= 12'h603;
      20'h05209: out <= 12'h603;
      20'h0520a: out <= 12'h603;
      20'h0520b: out <= 12'h603;
      20'h0520c: out <= 12'h222;
      20'h0520d: out <= 12'h222;
      20'h0520e: out <= 12'h222;
      20'h0520f: out <= 12'h222;
      20'h05210: out <= 12'h222;
      20'h05211: out <= 12'h222;
      20'h05212: out <= 12'h222;
      20'h05213: out <= 12'h222;
      20'h05214: out <= 12'h603;
      20'h05215: out <= 12'h603;
      20'h05216: out <= 12'h603;
      20'h05217: out <= 12'h603;
      20'h05218: out <= 12'h603;
      20'h05219: out <= 12'h603;
      20'h0521a: out <= 12'h603;
      20'h0521b: out <= 12'h603;
      20'h0521c: out <= 12'h000;
      20'h0521d: out <= 12'h000;
      20'h0521e: out <= 12'h000;
      20'h0521f: out <= 12'h6af;
      20'h05220: out <= 12'h6af;
      20'h05221: out <= 12'h000;
      20'h05222: out <= 12'h000;
      20'h05223: out <= 12'h000;
      20'h05224: out <= 12'h603;
      20'h05225: out <= 12'h603;
      20'h05226: out <= 12'h603;
      20'h05227: out <= 12'h603;
      20'h05228: out <= 12'h222;
      20'h05229: out <= 12'h222;
      20'h0522a: out <= 12'h222;
      20'h0522b: out <= 12'h222;
      20'h0522c: out <= 12'h222;
      20'h0522d: out <= 12'h222;
      20'h0522e: out <= 12'h222;
      20'h0522f: out <= 12'h222;
      20'h05230: out <= 12'h222;
      20'h05231: out <= 12'h222;
      20'h05232: out <= 12'h222;
      20'h05233: out <= 12'h222;
      20'h05234: out <= 12'h222;
      20'h05235: out <= 12'h222;
      20'h05236: out <= 12'h222;
      20'h05237: out <= 12'h222;
      20'h05238: out <= 12'h603;
      20'h05239: out <= 12'h603;
      20'h0523a: out <= 12'h603;
      20'h0523b: out <= 12'h603;
      20'h0523c: out <= 12'h000;
      20'h0523d: out <= 12'h000;
      20'h0523e: out <= 12'h000;
      20'h0523f: out <= 12'h16d;
      20'h05240: out <= 12'h16d;
      20'h05241: out <= 12'h16d;
      20'h05242: out <= 12'h000;
      20'h05243: out <= 12'h000;
      20'h05244: out <= 12'h603;
      20'h05245: out <= 12'h603;
      20'h05246: out <= 12'h603;
      20'h05247: out <= 12'h603;
      20'h05248: out <= 12'h222;
      20'h05249: out <= 12'h222;
      20'h0524a: out <= 12'h222;
      20'h0524b: out <= 12'h222;
      20'h0524c: out <= 12'h222;
      20'h0524d: out <= 12'h222;
      20'h0524e: out <= 12'h222;
      20'h0524f: out <= 12'h222;
      20'h05250: out <= 12'h222;
      20'h05251: out <= 12'h222;
      20'h05252: out <= 12'h222;
      20'h05253: out <= 12'h222;
      20'h05254: out <= 12'h222;
      20'h05255: out <= 12'h222;
      20'h05256: out <= 12'h222;
      20'h05257: out <= 12'h222;
      20'h05258: out <= 12'h603;
      20'h05259: out <= 12'h603;
      20'h0525a: out <= 12'h603;
      20'h0525b: out <= 12'h603;
      20'h0525c: out <= 12'h000;
      20'h0525d: out <= 12'h000;
      20'h0525e: out <= 12'h000;
      20'h0525f: out <= 12'h660;
      20'h05260: out <= 12'hbb0;
      20'h05261: out <= 12'h660;
      20'h05262: out <= 12'h000;
      20'h05263: out <= 12'h000;
      20'h05264: out <= 12'h603;
      20'h05265: out <= 12'h603;
      20'h05266: out <= 12'h603;
      20'h05267: out <= 12'h603;
      20'h05268: out <= 12'h222;
      20'h05269: out <= 12'h222;
      20'h0526a: out <= 12'h222;
      20'h0526b: out <= 12'h222;
      20'h0526c: out <= 12'h660;
      20'h0526d: out <= 12'h222;
      20'h0526e: out <= 12'h222;
      20'h0526f: out <= 12'h222;
      20'h05270: out <= 12'h222;
      20'h05271: out <= 12'h222;
      20'h05272: out <= 12'h222;
      20'h05273: out <= 12'h222;
      20'h05274: out <= 12'h660;
      20'h05275: out <= 12'h222;
      20'h05276: out <= 12'h222;
      20'h05277: out <= 12'h222;
      20'h05278: out <= 12'h000;
      20'h05279: out <= 12'h000;
      20'h0527a: out <= 12'h000;
      20'h0527b: out <= 12'h000;
      20'h0527c: out <= 12'h000;
      20'h0527d: out <= 12'h000;
      20'h0527e: out <= 12'h660;
      20'h0527f: out <= 12'hbb0;
      20'h05280: out <= 12'hee9;
      20'h05281: out <= 12'hbb0;
      20'h05282: out <= 12'h660;
      20'h05283: out <= 12'h000;
      20'h05284: out <= 12'h000;
      20'h05285: out <= 12'h000;
      20'h05286: out <= 12'h000;
      20'h05287: out <= 12'h000;
      20'h05288: out <= 12'h603;
      20'h05289: out <= 12'h603;
      20'h0528a: out <= 12'h603;
      20'h0528b: out <= 12'h603;
      20'h0528c: out <= 12'h000;
      20'h0528d: out <= 12'h666;
      20'h0528e: out <= 12'h666;
      20'h0528f: out <= 12'h666;
      20'h05290: out <= 12'h666;
      20'h05291: out <= 12'h666;
      20'h05292: out <= 12'h666;
      20'h05293: out <= 12'h666;
      20'h05294: out <= 12'h666;
      20'h05295: out <= 12'h666;
      20'h05296: out <= 12'h666;
      20'h05297: out <= 12'h666;
      20'h05298: out <= 12'h666;
      20'h05299: out <= 12'h666;
      20'h0529a: out <= 12'h666;
      20'h0529b: out <= 12'h666;
      20'h0529c: out <= 12'h000;
      20'h0529d: out <= 12'h000;
      20'h0529e: out <= 12'h000;
      20'h0529f: out <= 12'hb27;
      20'h052a0: out <= 12'hf87;
      20'h052a1: out <= 12'hee9;
      20'h052a2: out <= 12'hee9;
      20'h052a3: out <= 12'hf87;
      20'h052a4: out <= 12'hf87;
      20'h052a5: out <= 12'hf87;
      20'h052a6: out <= 12'hb27;
      20'h052a7: out <= 12'hb27;
      20'h052a8: out <= 12'hf87;
      20'h052a9: out <= 12'hee9;
      20'h052aa: out <= 12'h000;
      20'h052ab: out <= 12'h000;
      20'h052ac: out <= 12'h000;
      20'h052ad: out <= 12'h000;
      20'h052ae: out <= 12'h000;
      20'h052af: out <= 12'h000;
      20'h052b0: out <= 12'hb27;
      20'h052b1: out <= 12'hf87;
      20'h052b2: out <= 12'hf87;
      20'h052b3: out <= 12'hee9;
      20'h052b4: out <= 12'hee9;
      20'h052b5: out <= 12'hf87;
      20'h052b6: out <= 12'hf87;
      20'h052b7: out <= 12'hb27;
      20'h052b8: out <= 12'hb27;
      20'h052b9: out <= 12'hee9;
      20'h052ba: out <= 12'h000;
      20'h052bb: out <= 12'h000;
      20'h052bc: out <= 12'h603;
      20'h052bd: out <= 12'h603;
      20'h052be: out <= 12'h603;
      20'h052bf: out <= 12'h603;
      20'h052c0: out <= 12'h603;
      20'h052c1: out <= 12'h603;
      20'h052c2: out <= 12'h603;
      20'h052c3: out <= 12'h603;
      20'h052c4: out <= 12'h603;
      20'h052c5: out <= 12'h603;
      20'h052c6: out <= 12'h603;
      20'h052c7: out <= 12'h603;
      20'h052c8: out <= 12'h603;
      20'h052c9: out <= 12'h603;
      20'h052ca: out <= 12'h603;
      20'h052cb: out <= 12'h603;
      20'h052cc: out <= 12'h603;
      20'h052cd: out <= 12'h603;
      20'h052ce: out <= 12'h603;
      20'h052cf: out <= 12'h603;
      20'h052d0: out <= 12'h603;
      20'h052d1: out <= 12'h603;
      20'h052d2: out <= 12'h603;
      20'h052d3: out <= 12'h603;
      20'h052d4: out <= 12'h603;
      20'h052d5: out <= 12'h603;
      20'h052d6: out <= 12'h603;
      20'h052d7: out <= 12'h603;
      20'h052d8: out <= 12'h603;
      20'h052d9: out <= 12'h603;
      20'h052da: out <= 12'h603;
      20'h052db: out <= 12'h603;
      20'h052dc: out <= 12'h603;
      20'h052dd: out <= 12'h603;
      20'h052de: out <= 12'h603;
      20'h052df: out <= 12'h603;
      20'h052e0: out <= 12'hee9;
      20'h052e1: out <= 12'hf87;
      20'h052e2: out <= 12'hee9;
      20'h052e3: out <= 12'hf87;
      20'h052e4: out <= 12'hf87;
      20'h052e5: out <= 12'hb27;
      20'h052e6: out <= 12'hf87;
      20'h052e7: out <= 12'hb27;
      20'h052e8: out <= 12'h000;
      20'h052e9: out <= 12'h000;
      20'h052ea: out <= 12'h000;
      20'h052eb: out <= 12'h000;
      20'h052ec: out <= 12'h000;
      20'h052ed: out <= 12'h000;
      20'h052ee: out <= 12'h000;
      20'h052ef: out <= 12'h000;
      20'h052f0: out <= 12'h000;
      20'h052f1: out <= 12'h6af;
      20'h052f2: out <= 12'h16d;
      20'h052f3: out <= 12'h6af;
      20'h052f4: out <= 12'h000;
      20'h052f5: out <= 12'h000;
      20'h052f6: out <= 12'h000;
      20'h052f7: out <= 12'h16d;
      20'h052f8: out <= 12'hfff;
      20'h052f9: out <= 12'h16d;
      20'h052fa: out <= 12'h000;
      20'h052fb: out <= 12'h000;
      20'h052fc: out <= 12'h000;
      20'h052fd: out <= 12'h6af;
      20'h052fe: out <= 12'h16d;
      20'h052ff: out <= 12'h6af;
      20'h05300: out <= 12'h000;
      20'h05301: out <= 12'h000;
      20'h05302: out <= 12'h000;
      20'h05303: out <= 12'h000;
      20'h05304: out <= 12'h000;
      20'h05305: out <= 12'h000;
      20'h05306: out <= 12'h000;
      20'h05307: out <= 12'h000;
      20'h05308: out <= 12'h000;
      20'h05309: out <= 12'h000;
      20'h0530a: out <= 12'h000;
      20'h0530b: out <= 12'h000;
      20'h0530c: out <= 12'h000;
      20'h0530d: out <= 12'h000;
      20'h0530e: out <= 12'h000;
      20'h0530f: out <= 12'h000;
      20'h05310: out <= 12'h000;
      20'h05311: out <= 12'h000;
      20'h05312: out <= 12'h000;
      20'h05313: out <= 12'h000;
      20'h05314: out <= 12'h000;
      20'h05315: out <= 12'h000;
      20'h05316: out <= 12'h000;
      20'h05317: out <= 12'h000;
      20'h05318: out <= 12'h000;
      20'h05319: out <= 12'h000;
      20'h0531a: out <= 12'h000;
      20'h0531b: out <= 12'h000;
      20'h0531c: out <= 12'h000;
      20'h0531d: out <= 12'h000;
      20'h0531e: out <= 12'h000;
      20'h0531f: out <= 12'h000;
      20'h05320: out <= 12'h603;
      20'h05321: out <= 12'h603;
      20'h05322: out <= 12'h603;
      20'h05323: out <= 12'h603;
      20'h05324: out <= 12'h603;
      20'h05325: out <= 12'h603;
      20'h05326: out <= 12'h603;
      20'h05327: out <= 12'h603;
      20'h05328: out <= 12'h603;
      20'h05329: out <= 12'h603;
      20'h0532a: out <= 12'h603;
      20'h0532b: out <= 12'h603;
      20'h0532c: out <= 12'h603;
      20'h0532d: out <= 12'h603;
      20'h0532e: out <= 12'h603;
      20'h0532f: out <= 12'h603;
      20'h05330: out <= 12'h603;
      20'h05331: out <= 12'h603;
      20'h05332: out <= 12'h603;
      20'h05333: out <= 12'h603;
      20'h05334: out <= 12'h603;
      20'h05335: out <= 12'h603;
      20'h05336: out <= 12'h603;
      20'h05337: out <= 12'h603;
      20'h05338: out <= 12'h603;
      20'h05339: out <= 12'h603;
      20'h0533a: out <= 12'h603;
      20'h0533b: out <= 12'h603;
      20'h0533c: out <= 12'h603;
      20'h0533d: out <= 12'h603;
      20'h0533e: out <= 12'h603;
      20'h0533f: out <= 12'h603;
      20'h05340: out <= 12'h603;
      20'h05341: out <= 12'h603;
      20'h05342: out <= 12'h603;
      20'h05343: out <= 12'h603;
      20'h05344: out <= 12'h603;
      20'h05345: out <= 12'h603;
      20'h05346: out <= 12'h603;
      20'h05347: out <= 12'h603;
      20'h05348: out <= 12'h603;
      20'h05349: out <= 12'h603;
      20'h0534a: out <= 12'h603;
      20'h0534b: out <= 12'h603;
      20'h0534c: out <= 12'h603;
      20'h0534d: out <= 12'h603;
      20'h0534e: out <= 12'h603;
      20'h0534f: out <= 12'h603;
      20'h05350: out <= 12'h603;
      20'h05351: out <= 12'h603;
      20'h05352: out <= 12'h603;
      20'h05353: out <= 12'h603;
      20'h05354: out <= 12'h000;
      20'h05355: out <= 12'h000;
      20'h05356: out <= 12'h16d;
      20'h05357: out <= 12'h6af;
      20'h05358: out <= 12'hfff;
      20'h05359: out <= 12'h6af;
      20'h0535a: out <= 12'h16d;
      20'h0535b: out <= 12'h000;
      20'h0535c: out <= 12'h603;
      20'h0535d: out <= 12'h603;
      20'h0535e: out <= 12'h603;
      20'h0535f: out <= 12'h603;
      20'h05360: out <= 12'h603;
      20'h05361: out <= 12'h603;
      20'h05362: out <= 12'h603;
      20'h05363: out <= 12'h603;
      20'h05364: out <= 12'h603;
      20'h05365: out <= 12'h603;
      20'h05366: out <= 12'h603;
      20'h05367: out <= 12'h603;
      20'h05368: out <= 12'h603;
      20'h05369: out <= 12'h603;
      20'h0536a: out <= 12'h603;
      20'h0536b: out <= 12'h603;
      20'h0536c: out <= 12'h603;
      20'h0536d: out <= 12'h603;
      20'h0536e: out <= 12'h603;
      20'h0536f: out <= 12'h603;
      20'h05370: out <= 12'h603;
      20'h05371: out <= 12'h603;
      20'h05372: out <= 12'h603;
      20'h05373: out <= 12'h603;
      20'h05374: out <= 12'h000;
      20'h05375: out <= 12'h000;
      20'h05376: out <= 12'h000;
      20'h05377: out <= 12'h660;
      20'h05378: out <= 12'hbb0;
      20'h05379: out <= 12'h660;
      20'h0537a: out <= 12'h000;
      20'h0537b: out <= 12'h000;
      20'h0537c: out <= 12'h603;
      20'h0537d: out <= 12'h603;
      20'h0537e: out <= 12'h603;
      20'h0537f: out <= 12'h603;
      20'h05380: out <= 12'h222;
      20'h05381: out <= 12'h222;
      20'h05382: out <= 12'h222;
      20'h05383: out <= 12'h222;
      20'h05384: out <= 12'h222;
      20'h05385: out <= 12'h222;
      20'h05386: out <= 12'h222;
      20'h05387: out <= 12'h222;
      20'h05388: out <= 12'h222;
      20'h05389: out <= 12'h222;
      20'h0538a: out <= 12'h222;
      20'h0538b: out <= 12'h222;
      20'h0538c: out <= 12'h222;
      20'h0538d: out <= 12'h222;
      20'h0538e: out <= 12'h222;
      20'h0538f: out <= 12'h222;
      20'h05390: out <= 12'h000;
      20'h05391: out <= 12'h000;
      20'h05392: out <= 12'h000;
      20'h05393: out <= 12'h000;
      20'h05394: out <= 12'h000;
      20'h05395: out <= 12'h000;
      20'h05396: out <= 12'h000;
      20'h05397: out <= 12'h660;
      20'h05398: out <= 12'hee9;
      20'h05399: out <= 12'h660;
      20'h0539a: out <= 12'h000;
      20'h0539b: out <= 12'h000;
      20'h0539c: out <= 12'h000;
      20'h0539d: out <= 12'h000;
      20'h0539e: out <= 12'h000;
      20'h0539f: out <= 12'h000;
      20'h053a0: out <= 12'h603;
      20'h053a1: out <= 12'h603;
      20'h053a2: out <= 12'h603;
      20'h053a3: out <= 12'h603;
      20'h053a4: out <= 12'h000;
      20'h053a5: out <= 12'h000;
      20'h053a6: out <= 12'h000;
      20'h053a7: out <= 12'h000;
      20'h053a8: out <= 12'h000;
      20'h053a9: out <= 12'h000;
      20'h053aa: out <= 12'h666;
      20'h053ab: out <= 12'hbbb;
      20'h053ac: out <= 12'hfff;
      20'h053ad: out <= 12'hbbb;
      20'h053ae: out <= 12'h666;
      20'h053af: out <= 12'h000;
      20'h053b0: out <= 12'h000;
      20'h053b1: out <= 12'h000;
      20'h053b2: out <= 12'h000;
      20'h053b3: out <= 12'h000;
      20'h053b4: out <= 12'h000;
      20'h053b5: out <= 12'h000;
      20'h053b6: out <= 12'h000;
      20'h053b7: out <= 12'hb27;
      20'h053b8: out <= 12'hf87;
      20'h053b9: out <= 12'hee9;
      20'h053ba: out <= 12'hee9;
      20'h053bb: out <= 12'hf87;
      20'h053bc: out <= 12'hf87;
      20'h053bd: out <= 12'hf87;
      20'h053be: out <= 12'hb27;
      20'h053bf: out <= 12'hb27;
      20'h053c0: out <= 12'hf87;
      20'h053c1: out <= 12'hee9;
      20'h053c2: out <= 12'h000;
      20'h053c3: out <= 12'h000;
      20'h053c4: out <= 12'h000;
      20'h053c5: out <= 12'h000;
      20'h053c6: out <= 12'h000;
      20'h053c7: out <= 12'hb27;
      20'h053c8: out <= 12'hf87;
      20'h053c9: out <= 12'hf87;
      20'h053ca: out <= 12'hee9;
      20'h053cb: out <= 12'hee9;
      20'h053cc: out <= 12'hf87;
      20'h053cd: out <= 12'hf87;
      20'h053ce: out <= 12'hb27;
      20'h053cf: out <= 12'hb27;
      20'h053d0: out <= 12'hf87;
      20'h053d1: out <= 12'hee9;
      20'h053d2: out <= 12'h000;
      20'h053d3: out <= 12'h000;
      20'h053d4: out <= 12'h603;
      20'h053d5: out <= 12'h603;
      20'h053d6: out <= 12'h603;
      20'h053d7: out <= 12'h603;
      20'h053d8: out <= 12'h603;
      20'h053d9: out <= 12'h603;
      20'h053da: out <= 12'h603;
      20'h053db: out <= 12'h603;
      20'h053dc: out <= 12'h603;
      20'h053dd: out <= 12'h603;
      20'h053de: out <= 12'h603;
      20'h053df: out <= 12'h603;
      20'h053e0: out <= 12'h603;
      20'h053e1: out <= 12'h603;
      20'h053e2: out <= 12'h603;
      20'h053e3: out <= 12'h603;
      20'h053e4: out <= 12'h603;
      20'h053e5: out <= 12'h603;
      20'h053e6: out <= 12'h603;
      20'h053e7: out <= 12'h603;
      20'h053e8: out <= 12'h603;
      20'h053e9: out <= 12'h603;
      20'h053ea: out <= 12'h603;
      20'h053eb: out <= 12'h603;
      20'h053ec: out <= 12'h603;
      20'h053ed: out <= 12'h603;
      20'h053ee: out <= 12'h603;
      20'h053ef: out <= 12'h603;
      20'h053f0: out <= 12'h603;
      20'h053f1: out <= 12'h603;
      20'h053f2: out <= 12'h603;
      20'h053f3: out <= 12'h603;
      20'h053f4: out <= 12'h603;
      20'h053f5: out <= 12'h603;
      20'h053f6: out <= 12'h603;
      20'h053f7: out <= 12'h603;
      20'h053f8: out <= 12'hee9;
      20'h053f9: out <= 12'hf87;
      20'h053fa: out <= 12'hee9;
      20'h053fb: out <= 12'hf87;
      20'h053fc: out <= 12'hf87;
      20'h053fd: out <= 12'hb27;
      20'h053fe: out <= 12'hf87;
      20'h053ff: out <= 12'hb27;
      20'h05400: out <= 12'h000;
      20'h05401: out <= 12'h000;
      20'h05402: out <= 12'h000;
      20'h05403: out <= 12'h000;
      20'h05404: out <= 12'h000;
      20'h05405: out <= 12'h000;
      20'h05406: out <= 12'h000;
      20'h05407: out <= 12'h000;
      20'h05408: out <= 12'h000;
      20'h05409: out <= 12'h6af;
      20'h0540a: out <= 12'hfff;
      20'h0540b: out <= 12'h6af;
      20'h0540c: out <= 12'h000;
      20'h0540d: out <= 12'h16d;
      20'h0540e: out <= 12'h16d;
      20'h0540f: out <= 12'h16d;
      20'h05410: out <= 12'hfff;
      20'h05411: out <= 12'h16d;
      20'h05412: out <= 12'h16d;
      20'h05413: out <= 12'h16d;
      20'h05414: out <= 12'h000;
      20'h05415: out <= 12'h6af;
      20'h05416: out <= 12'hfff;
      20'h05417: out <= 12'h6af;
      20'h05418: out <= 12'h000;
      20'h05419: out <= 12'h000;
      20'h0541a: out <= 12'h000;
      20'h0541b: out <= 12'h000;
      20'h0541c: out <= 12'h000;
      20'h0541d: out <= 12'h000;
      20'h0541e: out <= 12'h000;
      20'h0541f: out <= 12'h000;
      20'h05420: out <= 12'h000;
      20'h05421: out <= 12'h000;
      20'h05422: out <= 12'h000;
      20'h05423: out <= 12'h000;
      20'h05424: out <= 12'h000;
      20'h05425: out <= 12'h000;
      20'h05426: out <= 12'h000;
      20'h05427: out <= 12'h000;
      20'h05428: out <= 12'h000;
      20'h05429: out <= 12'h000;
      20'h0542a: out <= 12'h000;
      20'h0542b: out <= 12'h000;
      20'h0542c: out <= 12'h000;
      20'h0542d: out <= 12'h000;
      20'h0542e: out <= 12'h000;
      20'h0542f: out <= 12'h000;
      20'h05430: out <= 12'h000;
      20'h05431: out <= 12'h000;
      20'h05432: out <= 12'h000;
      20'h05433: out <= 12'h000;
      20'h05434: out <= 12'h000;
      20'h05435: out <= 12'h000;
      20'h05436: out <= 12'h000;
      20'h05437: out <= 12'h000;
      20'h05438: out <= 12'h603;
      20'h05439: out <= 12'h603;
      20'h0543a: out <= 12'h603;
      20'h0543b: out <= 12'h603;
      20'h0543c: out <= 12'h603;
      20'h0543d: out <= 12'h603;
      20'h0543e: out <= 12'h603;
      20'h0543f: out <= 12'h603;
      20'h05440: out <= 12'h603;
      20'h05441: out <= 12'h603;
      20'h05442: out <= 12'h603;
      20'h05443: out <= 12'h603;
      20'h05444: out <= 12'h603;
      20'h05445: out <= 12'h603;
      20'h05446: out <= 12'h603;
      20'h05447: out <= 12'h603;
      20'h05448: out <= 12'h603;
      20'h05449: out <= 12'h603;
      20'h0544a: out <= 12'h603;
      20'h0544b: out <= 12'h603;
      20'h0544c: out <= 12'h603;
      20'h0544d: out <= 12'h603;
      20'h0544e: out <= 12'h603;
      20'h0544f: out <= 12'h603;
      20'h05450: out <= 12'h603;
      20'h05451: out <= 12'h603;
      20'h05452: out <= 12'h603;
      20'h05453: out <= 12'h603;
      20'h05454: out <= 12'h603;
      20'h05455: out <= 12'h603;
      20'h05456: out <= 12'h603;
      20'h05457: out <= 12'h603;
      20'h05458: out <= 12'h603;
      20'h05459: out <= 12'h603;
      20'h0545a: out <= 12'h603;
      20'h0545b: out <= 12'h603;
      20'h0545c: out <= 12'h603;
      20'h0545d: out <= 12'h603;
      20'h0545e: out <= 12'h603;
      20'h0545f: out <= 12'h603;
      20'h05460: out <= 12'h603;
      20'h05461: out <= 12'h603;
      20'h05462: out <= 12'h603;
      20'h05463: out <= 12'h603;
      20'h05464: out <= 12'h603;
      20'h05465: out <= 12'h603;
      20'h05466: out <= 12'h603;
      20'h05467: out <= 12'h603;
      20'h05468: out <= 12'h603;
      20'h05469: out <= 12'h603;
      20'h0546a: out <= 12'h603;
      20'h0546b: out <= 12'h603;
      20'h0546c: out <= 12'h000;
      20'h0546d: out <= 12'h6af;
      20'h0546e: out <= 12'h16d;
      20'h0546f: out <= 12'h6af;
      20'h05470: out <= 12'hfff;
      20'h05471: out <= 12'h6af;
      20'h05472: out <= 12'h16d;
      20'h05473: out <= 12'h6af;
      20'h05474: out <= 12'h603;
      20'h05475: out <= 12'h603;
      20'h05476: out <= 12'h603;
      20'h05477: out <= 12'h603;
      20'h05478: out <= 12'h603;
      20'h05479: out <= 12'h603;
      20'h0547a: out <= 12'h603;
      20'h0547b: out <= 12'h603;
      20'h0547c: out <= 12'h603;
      20'h0547d: out <= 12'h603;
      20'h0547e: out <= 12'h603;
      20'h0547f: out <= 12'h603;
      20'h05480: out <= 12'h603;
      20'h05481: out <= 12'h603;
      20'h05482: out <= 12'h603;
      20'h05483: out <= 12'h603;
      20'h05484: out <= 12'h603;
      20'h05485: out <= 12'h603;
      20'h05486: out <= 12'h603;
      20'h05487: out <= 12'h603;
      20'h05488: out <= 12'h603;
      20'h05489: out <= 12'h603;
      20'h0548a: out <= 12'h603;
      20'h0548b: out <= 12'h603;
      20'h0548c: out <= 12'h000;
      20'h0548d: out <= 12'h000;
      20'h0548e: out <= 12'h000;
      20'h0548f: out <= 12'h000;
      20'h05490: out <= 12'hbb0;
      20'h05491: out <= 12'h000;
      20'h05492: out <= 12'h000;
      20'h05493: out <= 12'h000;
      20'h05494: out <= 12'h603;
      20'h05495: out <= 12'h603;
      20'h05496: out <= 12'h603;
      20'h05497: out <= 12'h603;
      20'h05498: out <= 12'h222;
      20'h05499: out <= 12'h222;
      20'h0549a: out <= 12'h222;
      20'h0549b: out <= 12'h222;
      20'h0549c: out <= 12'h222;
      20'h0549d: out <= 12'h222;
      20'h0549e: out <= 12'h222;
      20'h0549f: out <= 12'h222;
      20'h054a0: out <= 12'h222;
      20'h054a1: out <= 12'h222;
      20'h054a2: out <= 12'h222;
      20'h054a3: out <= 12'h222;
      20'h054a4: out <= 12'h222;
      20'h054a5: out <= 12'h222;
      20'h054a6: out <= 12'h222;
      20'h054a7: out <= 12'h222;
      20'h054a8: out <= 12'h000;
      20'h054a9: out <= 12'h000;
      20'h054aa: out <= 12'h000;
      20'h054ab: out <= 12'h000;
      20'h054ac: out <= 12'h000;
      20'h054ad: out <= 12'h000;
      20'h054ae: out <= 12'h000;
      20'h054af: out <= 12'h000;
      20'h054b0: out <= 12'hbb0;
      20'h054b1: out <= 12'h000;
      20'h054b2: out <= 12'h000;
      20'h054b3: out <= 12'h000;
      20'h054b4: out <= 12'h000;
      20'h054b5: out <= 12'h000;
      20'h054b6: out <= 12'h000;
      20'h054b7: out <= 12'h000;
      20'h054b8: out <= 12'h603;
      20'h054b9: out <= 12'h603;
      20'h054ba: out <= 12'h603;
      20'h054bb: out <= 12'h603;
      20'h054bc: out <= 12'h000;
      20'h054bd: out <= 12'h000;
      20'h054be: out <= 12'h000;
      20'h054bf: out <= 12'h000;
      20'h054c0: out <= 12'h000;
      20'h054c1: out <= 12'h000;
      20'h054c2: out <= 12'h666;
      20'h054c3: out <= 12'hbbb;
      20'h054c4: out <= 12'hfff;
      20'h054c5: out <= 12'hbbb;
      20'h054c6: out <= 12'h666;
      20'h054c7: out <= 12'h000;
      20'h054c8: out <= 12'h000;
      20'h054c9: out <= 12'h000;
      20'h054ca: out <= 12'h000;
      20'h054cb: out <= 12'h000;
      20'h054cc: out <= 12'h000;
      20'h054cd: out <= 12'h000;
      20'h054ce: out <= 12'h000;
      20'h054cf: out <= 12'hb27;
      20'h054d0: out <= 12'hb27;
      20'h054d1: out <= 12'hb27;
      20'h054d2: out <= 12'hb27;
      20'h054d3: out <= 12'hb27;
      20'h054d4: out <= 12'hb27;
      20'h054d5: out <= 12'hb27;
      20'h054d6: out <= 12'hb27;
      20'h054d7: out <= 12'hb27;
      20'h054d8: out <= 12'hb27;
      20'h054d9: out <= 12'hb27;
      20'h054da: out <= 12'h000;
      20'h054db: out <= 12'h000;
      20'h054dc: out <= 12'h000;
      20'h054dd: out <= 12'h000;
      20'h054de: out <= 12'h000;
      20'h054df: out <= 12'hb27;
      20'h054e0: out <= 12'hb27;
      20'h054e1: out <= 12'hb27;
      20'h054e2: out <= 12'hb27;
      20'h054e3: out <= 12'hb27;
      20'h054e4: out <= 12'hb27;
      20'h054e5: out <= 12'hb27;
      20'h054e6: out <= 12'hb27;
      20'h054e7: out <= 12'hb27;
      20'h054e8: out <= 12'hb27;
      20'h054e9: out <= 12'hb27;
      20'h054ea: out <= 12'h000;
      20'h054eb: out <= 12'h000;
      20'h054ec: out <= 12'h603;
      20'h054ed: out <= 12'h603;
      20'h054ee: out <= 12'h603;
      20'h054ef: out <= 12'h603;
      20'h054f0: out <= 12'h603;
      20'h054f1: out <= 12'h603;
      20'h054f2: out <= 12'h603;
      20'h054f3: out <= 12'h603;
      20'h054f4: out <= 12'h603;
      20'h054f5: out <= 12'h603;
      20'h054f6: out <= 12'h603;
      20'h054f7: out <= 12'h603;
      20'h054f8: out <= 12'h603;
      20'h054f9: out <= 12'h603;
      20'h054fa: out <= 12'h603;
      20'h054fb: out <= 12'h603;
      20'h054fc: out <= 12'h603;
      20'h054fd: out <= 12'h603;
      20'h054fe: out <= 12'h603;
      20'h054ff: out <= 12'h603;
      20'h05500: out <= 12'h603;
      20'h05501: out <= 12'h603;
      20'h05502: out <= 12'h603;
      20'h05503: out <= 12'h603;
      20'h05504: out <= 12'h603;
      20'h05505: out <= 12'h603;
      20'h05506: out <= 12'h603;
      20'h05507: out <= 12'h603;
      20'h05508: out <= 12'h603;
      20'h05509: out <= 12'h603;
      20'h0550a: out <= 12'h603;
      20'h0550b: out <= 12'h603;
      20'h0550c: out <= 12'h603;
      20'h0550d: out <= 12'h603;
      20'h0550e: out <= 12'h603;
      20'h0550f: out <= 12'h603;
      20'h05510: out <= 12'hee9;
      20'h05511: out <= 12'hf87;
      20'h05512: out <= 12'hee9;
      20'h05513: out <= 12'hb27;
      20'h05514: out <= 12'hb27;
      20'h05515: out <= 12'hb27;
      20'h05516: out <= 12'hf87;
      20'h05517: out <= 12'hb27;
      20'h05518: out <= 12'h000;
      20'h05519: out <= 12'h000;
      20'h0551a: out <= 12'h000;
      20'h0551b: out <= 12'h000;
      20'h0551c: out <= 12'h000;
      20'h0551d: out <= 12'h000;
      20'h0551e: out <= 12'h000;
      20'h0551f: out <= 12'h000;
      20'h05520: out <= 12'h000;
      20'h05521: out <= 12'h6af;
      20'h05522: out <= 12'h16d;
      20'h05523: out <= 12'h16d;
      20'h05524: out <= 12'h16d;
      20'h05525: out <= 12'hfff;
      20'h05526: out <= 12'h6af;
      20'h05527: out <= 12'h16d;
      20'h05528: out <= 12'h16d;
      20'h05529: out <= 12'h16d;
      20'h0552a: out <= 12'h6af;
      20'h0552b: out <= 12'hfff;
      20'h0552c: out <= 12'h16d;
      20'h0552d: out <= 12'h16d;
      20'h0552e: out <= 12'h16d;
      20'h0552f: out <= 12'h6af;
      20'h05530: out <= 12'h000;
      20'h05531: out <= 12'h000;
      20'h05532: out <= 12'h000;
      20'h05533: out <= 12'h000;
      20'h05534: out <= 12'h000;
      20'h05535: out <= 12'h000;
      20'h05536: out <= 12'h000;
      20'h05537: out <= 12'h000;
      20'h05538: out <= 12'h000;
      20'h05539: out <= 12'h000;
      20'h0553a: out <= 12'h000;
      20'h0553b: out <= 12'h000;
      20'h0553c: out <= 12'h000;
      20'h0553d: out <= 12'h000;
      20'h0553e: out <= 12'h000;
      20'h0553f: out <= 12'h000;
      20'h05540: out <= 12'h000;
      20'h05541: out <= 12'h000;
      20'h05542: out <= 12'h000;
      20'h05543: out <= 12'h000;
      20'h05544: out <= 12'h000;
      20'h05545: out <= 12'h000;
      20'h05546: out <= 12'h000;
      20'h05547: out <= 12'h000;
      20'h05548: out <= 12'h000;
      20'h05549: out <= 12'h000;
      20'h0554a: out <= 12'h000;
      20'h0554b: out <= 12'h000;
      20'h0554c: out <= 12'h000;
      20'h0554d: out <= 12'h000;
      20'h0554e: out <= 12'h000;
      20'h0554f: out <= 12'h000;
      20'h05550: out <= 12'h603;
      20'h05551: out <= 12'h603;
      20'h05552: out <= 12'h603;
      20'h05553: out <= 12'h603;
      20'h05554: out <= 12'h603;
      20'h05555: out <= 12'h603;
      20'h05556: out <= 12'h603;
      20'h05557: out <= 12'h603;
      20'h05558: out <= 12'h603;
      20'h05559: out <= 12'h603;
      20'h0555a: out <= 12'h603;
      20'h0555b: out <= 12'h603;
      20'h0555c: out <= 12'h603;
      20'h0555d: out <= 12'h603;
      20'h0555e: out <= 12'h603;
      20'h0555f: out <= 12'h603;
      20'h05560: out <= 12'h603;
      20'h05561: out <= 12'h603;
      20'h05562: out <= 12'h603;
      20'h05563: out <= 12'h603;
      20'h05564: out <= 12'h603;
      20'h05565: out <= 12'h603;
      20'h05566: out <= 12'h603;
      20'h05567: out <= 12'h603;
      20'h05568: out <= 12'h603;
      20'h05569: out <= 12'h603;
      20'h0556a: out <= 12'h603;
      20'h0556b: out <= 12'h603;
      20'h0556c: out <= 12'h603;
      20'h0556d: out <= 12'h603;
      20'h0556e: out <= 12'h603;
      20'h0556f: out <= 12'h603;
      20'h05570: out <= 12'h603;
      20'h05571: out <= 12'h603;
      20'h05572: out <= 12'h603;
      20'h05573: out <= 12'h603;
      20'h05574: out <= 12'h603;
      20'h05575: out <= 12'h603;
      20'h05576: out <= 12'h603;
      20'h05577: out <= 12'h603;
      20'h05578: out <= 12'h603;
      20'h05579: out <= 12'h603;
      20'h0557a: out <= 12'h603;
      20'h0557b: out <= 12'h603;
      20'h0557c: out <= 12'h603;
      20'h0557d: out <= 12'h603;
      20'h0557e: out <= 12'h603;
      20'h0557f: out <= 12'h603;
      20'h05580: out <= 12'h603;
      20'h05581: out <= 12'h603;
      20'h05582: out <= 12'h603;
      20'h05583: out <= 12'h603;
      20'h05584: out <= 12'h000;
      20'h05585: out <= 12'h6af;
      20'h05586: out <= 12'h16d;
      20'h05587: out <= 12'h6af;
      20'h05588: out <= 12'hfff;
      20'h05589: out <= 12'h6af;
      20'h0558a: out <= 12'h16d;
      20'h0558b: out <= 12'h6af;
      20'h0558c: out <= 12'h603;
      20'h0558d: out <= 12'h603;
      20'h0558e: out <= 12'h603;
      20'h0558f: out <= 12'h603;
      20'h05590: out <= 12'h603;
      20'h05591: out <= 12'h603;
      20'h05592: out <= 12'h603;
      20'h05593: out <= 12'h603;
      20'h05594: out <= 12'h603;
      20'h05595: out <= 12'h603;
      20'h05596: out <= 12'h603;
      20'h05597: out <= 12'h603;
      20'h05598: out <= 12'h603;
      20'h05599: out <= 12'h603;
      20'h0559a: out <= 12'h603;
      20'h0559b: out <= 12'h603;
      20'h0559c: out <= 12'h603;
      20'h0559d: out <= 12'h603;
      20'h0559e: out <= 12'h603;
      20'h0559f: out <= 12'h603;
      20'h055a0: out <= 12'h603;
      20'h055a1: out <= 12'h603;
      20'h055a2: out <= 12'h603;
      20'h055a3: out <= 12'h603;
      20'h055a4: out <= 12'h000;
      20'h055a5: out <= 12'h000;
      20'h055a6: out <= 12'h000;
      20'h055a7: out <= 12'h000;
      20'h055a8: out <= 12'h660;
      20'h055a9: out <= 12'h000;
      20'h055aa: out <= 12'h000;
      20'h055ab: out <= 12'h000;
      20'h055ac: out <= 12'h603;
      20'h055ad: out <= 12'h603;
      20'h055ae: out <= 12'h603;
      20'h055af: out <= 12'h603;
      20'h055b0: out <= 12'h222;
      20'h055b1: out <= 12'h222;
      20'h055b2: out <= 12'h222;
      20'h055b3: out <= 12'h222;
      20'h055b4: out <= 12'h222;
      20'h055b5: out <= 12'h222;
      20'h055b6: out <= 12'h222;
      20'h055b7: out <= 12'h222;
      20'h055b8: out <= 12'h222;
      20'h055b9: out <= 12'h222;
      20'h055ba: out <= 12'h222;
      20'h055bb: out <= 12'h222;
      20'h055bc: out <= 12'h222;
      20'h055bd: out <= 12'h222;
      20'h055be: out <= 12'h222;
      20'h055bf: out <= 12'h222;
      20'h055c0: out <= 12'h000;
      20'h055c1: out <= 12'h000;
      20'h055c2: out <= 12'h000;
      20'h055c3: out <= 12'h000;
      20'h055c4: out <= 12'h000;
      20'h055c5: out <= 12'h000;
      20'h055c6: out <= 12'h000;
      20'h055c7: out <= 12'h000;
      20'h055c8: out <= 12'h660;
      20'h055c9: out <= 12'h000;
      20'h055ca: out <= 12'h000;
      20'h055cb: out <= 12'h000;
      20'h055cc: out <= 12'h000;
      20'h055cd: out <= 12'h000;
      20'h055ce: out <= 12'h000;
      20'h055cf: out <= 12'h000;
      20'h055d0: out <= 12'h603;
      20'h055d1: out <= 12'h603;
      20'h055d2: out <= 12'h603;
      20'h055d3: out <= 12'h603;
      20'h055d4: out <= 12'h000;
      20'h055d5: out <= 12'h000;
      20'h055d6: out <= 12'h000;
      20'h055d7: out <= 12'h666;
      20'h055d8: out <= 12'h666;
      20'h055d9: out <= 12'hbbb;
      20'h055da: out <= 12'hbbb;
      20'h055db: out <= 12'hfff;
      20'h055dc: out <= 12'hfff;
      20'h055dd: out <= 12'hfff;
      20'h055de: out <= 12'hbbb;
      20'h055df: out <= 12'hbbb;
      20'h055e0: out <= 12'h666;
      20'h055e1: out <= 12'h666;
      20'h055e2: out <= 12'h000;
      20'h055e3: out <= 12'h000;
      20'h055e4: out <= 12'h000;
      20'h055e5: out <= 12'h000;
      20'h055e6: out <= 12'hb27;
      20'h055e7: out <= 12'hf87;
      20'h055e8: out <= 12'hee9;
      20'h055e9: out <= 12'hee9;
      20'h055ea: out <= 12'hf87;
      20'h055eb: out <= 12'hf87;
      20'h055ec: out <= 12'hf87;
      20'h055ed: out <= 12'hf87;
      20'h055ee: out <= 12'hf87;
      20'h055ef: out <= 12'hb27;
      20'h055f0: out <= 12'hb27;
      20'h055f1: out <= 12'hf87;
      20'h055f2: out <= 12'hee9;
      20'h055f3: out <= 12'h000;
      20'h055f4: out <= 12'h000;
      20'h055f5: out <= 12'h000;
      20'h055f6: out <= 12'hb27;
      20'h055f7: out <= 12'hf87;
      20'h055f8: out <= 12'hee9;
      20'h055f9: out <= 12'hee9;
      20'h055fa: out <= 12'hf87;
      20'h055fb: out <= 12'hf87;
      20'h055fc: out <= 12'hf87;
      20'h055fd: out <= 12'hf87;
      20'h055fe: out <= 12'hf87;
      20'h055ff: out <= 12'hb27;
      20'h05600: out <= 12'hb27;
      20'h05601: out <= 12'hf87;
      20'h05602: out <= 12'hee9;
      20'h05603: out <= 12'h000;
      20'h05604: out <= 12'h603;
      20'h05605: out <= 12'h603;
      20'h05606: out <= 12'h603;
      20'h05607: out <= 12'h603;
      20'h05608: out <= 12'h603;
      20'h05609: out <= 12'h603;
      20'h0560a: out <= 12'h603;
      20'h0560b: out <= 12'h603;
      20'h0560c: out <= 12'h603;
      20'h0560d: out <= 12'h603;
      20'h0560e: out <= 12'h603;
      20'h0560f: out <= 12'h603;
      20'h05610: out <= 12'h603;
      20'h05611: out <= 12'h603;
      20'h05612: out <= 12'h603;
      20'h05613: out <= 12'h603;
      20'h05614: out <= 12'h603;
      20'h05615: out <= 12'h603;
      20'h05616: out <= 12'h603;
      20'h05617: out <= 12'h603;
      20'h05618: out <= 12'h603;
      20'h05619: out <= 12'h603;
      20'h0561a: out <= 12'h603;
      20'h0561b: out <= 12'h603;
      20'h0561c: out <= 12'h603;
      20'h0561d: out <= 12'h603;
      20'h0561e: out <= 12'h603;
      20'h0561f: out <= 12'h603;
      20'h05620: out <= 12'h603;
      20'h05621: out <= 12'h603;
      20'h05622: out <= 12'h603;
      20'h05623: out <= 12'h603;
      20'h05624: out <= 12'h603;
      20'h05625: out <= 12'h603;
      20'h05626: out <= 12'h603;
      20'h05627: out <= 12'h603;
      20'h05628: out <= 12'hee9;
      20'h05629: out <= 12'hf87;
      20'h0562a: out <= 12'hf87;
      20'h0562b: out <= 12'hf87;
      20'h0562c: out <= 12'hf87;
      20'h0562d: out <= 12'hf87;
      20'h0562e: out <= 12'hf87;
      20'h0562f: out <= 12'hb27;
      20'h05630: out <= 12'h000;
      20'h05631: out <= 12'h000;
      20'h05632: out <= 12'h000;
      20'h05633: out <= 12'h000;
      20'h05634: out <= 12'h000;
      20'h05635: out <= 12'h000;
      20'h05636: out <= 12'h000;
      20'h05637: out <= 12'h000;
      20'h05638: out <= 12'h000;
      20'h05639: out <= 12'h6af;
      20'h0563a: out <= 12'hfff;
      20'h0563b: out <= 12'h16d;
      20'h0563c: out <= 12'hfff;
      20'h0563d: out <= 12'h6af;
      20'h0563e: out <= 12'h16d;
      20'h0563f: out <= 12'h16d;
      20'h05640: out <= 12'h6af;
      20'h05641: out <= 12'h16d;
      20'h05642: out <= 12'h16d;
      20'h05643: out <= 12'h6af;
      20'h05644: out <= 12'hfff;
      20'h05645: out <= 12'h16d;
      20'h05646: out <= 12'hfff;
      20'h05647: out <= 12'h6af;
      20'h05648: out <= 12'h000;
      20'h05649: out <= 12'h000;
      20'h0564a: out <= 12'h000;
      20'h0564b: out <= 12'h000;
      20'h0564c: out <= 12'h000;
      20'h0564d: out <= 12'h000;
      20'h0564e: out <= 12'h000;
      20'h0564f: out <= 12'h000;
      20'h05650: out <= 12'h000;
      20'h05651: out <= 12'h000;
      20'h05652: out <= 12'h000;
      20'h05653: out <= 12'h000;
      20'h05654: out <= 12'h000;
      20'h05655: out <= 12'h000;
      20'h05656: out <= 12'h000;
      20'h05657: out <= 12'h000;
      20'h05658: out <= 12'h000;
      20'h05659: out <= 12'h000;
      20'h0565a: out <= 12'h000;
      20'h0565b: out <= 12'h000;
      20'h0565c: out <= 12'h000;
      20'h0565d: out <= 12'h000;
      20'h0565e: out <= 12'h000;
      20'h0565f: out <= 12'h000;
      20'h05660: out <= 12'h000;
      20'h05661: out <= 12'h000;
      20'h05662: out <= 12'h000;
      20'h05663: out <= 12'h000;
      20'h05664: out <= 12'h000;
      20'h05665: out <= 12'h000;
      20'h05666: out <= 12'h000;
      20'h05667: out <= 12'h000;
      20'h05668: out <= 12'h603;
      20'h05669: out <= 12'h603;
      20'h0566a: out <= 12'h603;
      20'h0566b: out <= 12'h603;
      20'h0566c: out <= 12'h603;
      20'h0566d: out <= 12'h603;
      20'h0566e: out <= 12'h603;
      20'h0566f: out <= 12'h603;
      20'h05670: out <= 12'h603;
      20'h05671: out <= 12'h603;
      20'h05672: out <= 12'h603;
      20'h05673: out <= 12'h603;
      20'h05674: out <= 12'h603;
      20'h05675: out <= 12'h603;
      20'h05676: out <= 12'h603;
      20'h05677: out <= 12'h603;
      20'h05678: out <= 12'h603;
      20'h05679: out <= 12'h603;
      20'h0567a: out <= 12'h603;
      20'h0567b: out <= 12'h603;
      20'h0567c: out <= 12'h603;
      20'h0567d: out <= 12'h603;
      20'h0567e: out <= 12'h603;
      20'h0567f: out <= 12'h603;
      20'h05680: out <= 12'h603;
      20'h05681: out <= 12'h603;
      20'h05682: out <= 12'h603;
      20'h05683: out <= 12'h603;
      20'h05684: out <= 12'h603;
      20'h05685: out <= 12'h603;
      20'h05686: out <= 12'h603;
      20'h05687: out <= 12'h603;
      20'h05688: out <= 12'h603;
      20'h05689: out <= 12'h603;
      20'h0568a: out <= 12'h603;
      20'h0568b: out <= 12'h603;
      20'h0568c: out <= 12'h603;
      20'h0568d: out <= 12'h603;
      20'h0568e: out <= 12'h603;
      20'h0568f: out <= 12'h603;
      20'h05690: out <= 12'h603;
      20'h05691: out <= 12'h603;
      20'h05692: out <= 12'h603;
      20'h05693: out <= 12'h603;
      20'h05694: out <= 12'h603;
      20'h05695: out <= 12'h603;
      20'h05696: out <= 12'h603;
      20'h05697: out <= 12'h603;
      20'h05698: out <= 12'h603;
      20'h05699: out <= 12'h603;
      20'h0569a: out <= 12'h603;
      20'h0569b: out <= 12'h603;
      20'h0569c: out <= 12'h000;
      20'h0569d: out <= 12'h000;
      20'h0569e: out <= 12'h000;
      20'h0569f: out <= 12'h000;
      20'h056a0: out <= 12'h000;
      20'h056a1: out <= 12'h000;
      20'h056a2: out <= 12'h000;
      20'h056a3: out <= 12'h000;
      20'h056a4: out <= 12'h603;
      20'h056a5: out <= 12'h603;
      20'h056a6: out <= 12'h603;
      20'h056a7: out <= 12'h603;
      20'h056a8: out <= 12'h603;
      20'h056a9: out <= 12'h603;
      20'h056aa: out <= 12'h603;
      20'h056ab: out <= 12'h603;
      20'h056ac: out <= 12'h603;
      20'h056ad: out <= 12'h603;
      20'h056ae: out <= 12'h603;
      20'h056af: out <= 12'h603;
      20'h056b0: out <= 12'h603;
      20'h056b1: out <= 12'h603;
      20'h056b2: out <= 12'h603;
      20'h056b3: out <= 12'h603;
      20'h056b4: out <= 12'h603;
      20'h056b5: out <= 12'h603;
      20'h056b6: out <= 12'h603;
      20'h056b7: out <= 12'h603;
      20'h056b8: out <= 12'h603;
      20'h056b9: out <= 12'h603;
      20'h056ba: out <= 12'h603;
      20'h056bb: out <= 12'h603;
      20'h056bc: out <= 12'h000;
      20'h056bd: out <= 12'h000;
      20'h056be: out <= 12'h000;
      20'h056bf: out <= 12'h000;
      20'h056c0: out <= 12'h660;
      20'h056c1: out <= 12'h000;
      20'h056c2: out <= 12'h000;
      20'h056c3: out <= 12'h000;
      20'h056c4: out <= 12'h603;
      20'h056c5: out <= 12'h603;
      20'h056c6: out <= 12'h603;
      20'h056c7: out <= 12'h603;
      20'h056c8: out <= 12'h222;
      20'h056c9: out <= 12'h222;
      20'h056ca: out <= 12'h222;
      20'h056cb: out <= 12'h222;
      20'h056cc: out <= 12'h222;
      20'h056cd: out <= 12'h222;
      20'h056ce: out <= 12'h222;
      20'h056cf: out <= 12'h222;
      20'h056d0: out <= 12'h222;
      20'h056d1: out <= 12'h222;
      20'h056d2: out <= 12'h222;
      20'h056d3: out <= 12'h222;
      20'h056d4: out <= 12'h222;
      20'h056d5: out <= 12'h222;
      20'h056d6: out <= 12'h222;
      20'h056d7: out <= 12'h222;
      20'h056d8: out <= 12'h000;
      20'h056d9: out <= 12'h000;
      20'h056da: out <= 12'h000;
      20'h056db: out <= 12'h000;
      20'h056dc: out <= 12'h000;
      20'h056dd: out <= 12'h000;
      20'h056de: out <= 12'h000;
      20'h056df: out <= 12'h000;
      20'h056e0: out <= 12'h000;
      20'h056e1: out <= 12'h000;
      20'h056e2: out <= 12'h000;
      20'h056e3: out <= 12'h000;
      20'h056e4: out <= 12'h000;
      20'h056e5: out <= 12'h000;
      20'h056e6: out <= 12'h000;
      20'h056e7: out <= 12'h000;
      20'h056e8: out <= 12'h603;
      20'h056e9: out <= 12'h603;
      20'h056ea: out <= 12'h603;
      20'h056eb: out <= 12'h603;
      20'h056ec: out <= 12'h000;
      20'h056ed: out <= 12'h000;
      20'h056ee: out <= 12'h000;
      20'h056ef: out <= 12'h000;
      20'h056f0: out <= 12'h000;
      20'h056f1: out <= 12'h000;
      20'h056f2: out <= 12'h000;
      20'h056f3: out <= 12'h000;
      20'h056f4: out <= 12'h000;
      20'h056f5: out <= 12'h000;
      20'h056f6: out <= 12'h000;
      20'h056f7: out <= 12'h000;
      20'h056f8: out <= 12'h000;
      20'h056f9: out <= 12'h000;
      20'h056fa: out <= 12'h000;
      20'h056fb: out <= 12'h000;
      20'h056fc: out <= 12'h000;
      20'h056fd: out <= 12'h000;
      20'h056fe: out <= 12'h000;
      20'h056ff: out <= 12'h000;
      20'h05700: out <= 12'h000;
      20'h05701: out <= 12'h000;
      20'h05702: out <= 12'h000;
      20'h05703: out <= 12'h000;
      20'h05704: out <= 12'h000;
      20'h05705: out <= 12'h000;
      20'h05706: out <= 12'h000;
      20'h05707: out <= 12'h000;
      20'h05708: out <= 12'h000;
      20'h05709: out <= 12'h000;
      20'h0570a: out <= 12'h000;
      20'h0570b: out <= 12'h000;
      20'h0570c: out <= 12'h000;
      20'h0570d: out <= 12'h000;
      20'h0570e: out <= 12'h000;
      20'h0570f: out <= 12'h000;
      20'h05710: out <= 12'h000;
      20'h05711: out <= 12'h000;
      20'h05712: out <= 12'h000;
      20'h05713: out <= 12'h000;
      20'h05714: out <= 12'h000;
      20'h05715: out <= 12'h000;
      20'h05716: out <= 12'h000;
      20'h05717: out <= 12'h000;
      20'h05718: out <= 12'h000;
      20'h05719: out <= 12'h000;
      20'h0571a: out <= 12'h000;
      20'h0571b: out <= 12'h000;
      20'h0571c: out <= 12'h603;
      20'h0571d: out <= 12'h603;
      20'h0571e: out <= 12'h603;
      20'h0571f: out <= 12'h603;
      20'h05720: out <= 12'h603;
      20'h05721: out <= 12'h603;
      20'h05722: out <= 12'h603;
      20'h05723: out <= 12'h603;
      20'h05724: out <= 12'h603;
      20'h05725: out <= 12'h603;
      20'h05726: out <= 12'h603;
      20'h05727: out <= 12'h603;
      20'h05728: out <= 12'h603;
      20'h05729: out <= 12'h603;
      20'h0572a: out <= 12'h603;
      20'h0572b: out <= 12'h603;
      20'h0572c: out <= 12'h603;
      20'h0572d: out <= 12'h603;
      20'h0572e: out <= 12'h603;
      20'h0572f: out <= 12'h603;
      20'h05730: out <= 12'h603;
      20'h05731: out <= 12'h603;
      20'h05732: out <= 12'h603;
      20'h05733: out <= 12'h603;
      20'h05734: out <= 12'h603;
      20'h05735: out <= 12'h603;
      20'h05736: out <= 12'h603;
      20'h05737: out <= 12'h603;
      20'h05738: out <= 12'h603;
      20'h05739: out <= 12'h603;
      20'h0573a: out <= 12'h603;
      20'h0573b: out <= 12'h603;
      20'h0573c: out <= 12'h603;
      20'h0573d: out <= 12'h603;
      20'h0573e: out <= 12'h603;
      20'h0573f: out <= 12'h603;
      20'h05740: out <= 12'hb27;
      20'h05741: out <= 12'hb27;
      20'h05742: out <= 12'hb27;
      20'h05743: out <= 12'hb27;
      20'h05744: out <= 12'hb27;
      20'h05745: out <= 12'hb27;
      20'h05746: out <= 12'hb27;
      20'h05747: out <= 12'hb27;
      20'h05748: out <= 12'h000;
      20'h05749: out <= 12'h000;
      20'h0574a: out <= 12'h000;
      20'h0574b: out <= 12'h000;
      20'h0574c: out <= 12'h000;
      20'h0574d: out <= 12'h000;
      20'h0574e: out <= 12'h000;
      20'h0574f: out <= 12'h000;
      20'h05750: out <= 12'h000;
      20'h05751: out <= 12'h6af;
      20'h05752: out <= 12'h16d;
      20'h05753: out <= 12'h16d;
      20'h05754: out <= 12'h6af;
      20'h05755: out <= 12'h16d;
      20'h05756: out <= 12'h16d;
      20'h05757: out <= 12'h6af;
      20'h05758: out <= 12'hfff;
      20'h05759: out <= 12'h6af;
      20'h0575a: out <= 12'h16d;
      20'h0575b: out <= 12'h16d;
      20'h0575c: out <= 12'h6af;
      20'h0575d: out <= 12'h16d;
      20'h0575e: out <= 12'h16d;
      20'h0575f: out <= 12'h6af;
      20'h05760: out <= 12'h000;
      20'h05761: out <= 12'h000;
      20'h05762: out <= 12'h000;
      20'h05763: out <= 12'h000;
      20'h05764: out <= 12'h000;
      20'h05765: out <= 12'h000;
      20'h05766: out <= 12'h000;
      20'h05767: out <= 12'h000;
      20'h05768: out <= 12'h000;
      20'h05769: out <= 12'h000;
      20'h0576a: out <= 12'h000;
      20'h0576b: out <= 12'h000;
      20'h0576c: out <= 12'h000;
      20'h0576d: out <= 12'h000;
      20'h0576e: out <= 12'h000;
      20'h0576f: out <= 12'h000;
      20'h05770: out <= 12'h000;
      20'h05771: out <= 12'h000;
      20'h05772: out <= 12'h000;
      20'h05773: out <= 12'h000;
      20'h05774: out <= 12'h000;
      20'h05775: out <= 12'h000;
      20'h05776: out <= 12'h000;
      20'h05777: out <= 12'h000;
      20'h05778: out <= 12'h000;
      20'h05779: out <= 12'h000;
      20'h0577a: out <= 12'h000;
      20'h0577b: out <= 12'h000;
      20'h0577c: out <= 12'h000;
      20'h0577d: out <= 12'h000;
      20'h0577e: out <= 12'h000;
      20'h0577f: out <= 12'h000;
      20'h05780: out <= 12'h000;
      20'h05781: out <= 12'h000;
      20'h05782: out <= 12'h000;
      20'h05783: out <= 12'h000;
      20'h05784: out <= 12'h000;
      20'h05785: out <= 12'h000;
      20'h05786: out <= 12'h000;
      20'h05787: out <= 12'h000;
      20'h05788: out <= 12'h000;
      20'h05789: out <= 12'h000;
      20'h0578a: out <= 12'h000;
      20'h0578b: out <= 12'h000;
      20'h0578c: out <= 12'h000;
      20'h0578d: out <= 12'h000;
      20'h0578e: out <= 12'h000;
      20'h0578f: out <= 12'h000;
      20'h05790: out <= 12'h222;
      20'h05791: out <= 12'h222;
      20'h05792: out <= 12'h222;
      20'h05793: out <= 12'h222;
      20'h05794: out <= 12'h222;
      20'h05795: out <= 12'h222;
      20'h05796: out <= 12'h222;
      20'h05797: out <= 12'h222;
      20'h05798: out <= 12'h222;
      20'h05799: out <= 12'h222;
      20'h0579a: out <= 12'h222;
      20'h0579b: out <= 12'h222;
      20'h0579c: out <= 12'h222;
      20'h0579d: out <= 12'h222;
      20'h0579e: out <= 12'h222;
      20'h0579f: out <= 12'h222;
      20'h057a0: out <= 12'h000;
      20'h057a1: out <= 12'h000;
      20'h057a2: out <= 12'h000;
      20'h057a3: out <= 12'h000;
      20'h057a4: out <= 12'h000;
      20'h057a5: out <= 12'h000;
      20'h057a6: out <= 12'h000;
      20'h057a7: out <= 12'h666;
      20'h057a8: out <= 12'hfff;
      20'h057a9: out <= 12'h666;
      20'h057aa: out <= 12'h000;
      20'h057ab: out <= 12'h000;
      20'h057ac: out <= 12'h000;
      20'h057ad: out <= 12'h000;
      20'h057ae: out <= 12'h000;
      20'h057af: out <= 12'h000;
      20'h057b0: out <= 12'h222;
      20'h057b1: out <= 12'h222;
      20'h057b2: out <= 12'h222;
      20'h057b3: out <= 12'h222;
      20'h057b4: out <= 12'h222;
      20'h057b5: out <= 12'h222;
      20'h057b6: out <= 12'h222;
      20'h057b7: out <= 12'h666;
      20'h057b8: out <= 12'hfff;
      20'h057b9: out <= 12'h666;
      20'h057ba: out <= 12'h222;
      20'h057bb: out <= 12'h222;
      20'h057bc: out <= 12'h222;
      20'h057bd: out <= 12'h222;
      20'h057be: out <= 12'h222;
      20'h057bf: out <= 12'h222;
      20'h057c0: out <= 12'h000;
      20'h057c1: out <= 12'h000;
      20'h057c2: out <= 12'h000;
      20'h057c3: out <= 12'h000;
      20'h057c4: out <= 12'h000;
      20'h057c5: out <= 12'h000;
      20'h057c6: out <= 12'h000;
      20'h057c7: out <= 12'h000;
      20'h057c8: out <= 12'h000;
      20'h057c9: out <= 12'h000;
      20'h057ca: out <= 12'h000;
      20'h057cb: out <= 12'h000;
      20'h057cc: out <= 12'h000;
      20'h057cd: out <= 12'h000;
      20'h057ce: out <= 12'h000;
      20'h057cf: out <= 12'h000;
      20'h057d0: out <= 12'h222;
      20'h057d1: out <= 12'h222;
      20'h057d2: out <= 12'h222;
      20'h057d3: out <= 12'h222;
      20'h057d4: out <= 12'h222;
      20'h057d5: out <= 12'h222;
      20'h057d6: out <= 12'h222;
      20'h057d7: out <= 12'h222;
      20'h057d8: out <= 12'h222;
      20'h057d9: out <= 12'h222;
      20'h057da: out <= 12'h222;
      20'h057db: out <= 12'h222;
      20'h057dc: out <= 12'h222;
      20'h057dd: out <= 12'h222;
      20'h057de: out <= 12'h222;
      20'h057df: out <= 12'h222;
      20'h057e0: out <= 12'h000;
      20'h057e1: out <= 12'h000;
      20'h057e2: out <= 12'h000;
      20'h057e3: out <= 12'h000;
      20'h057e4: out <= 12'h000;
      20'h057e5: out <= 12'h000;
      20'h057e6: out <= 12'h000;
      20'h057e7: out <= 12'h000;
      20'h057e8: out <= 12'h000;
      20'h057e9: out <= 12'h000;
      20'h057ea: out <= 12'h000;
      20'h057eb: out <= 12'h000;
      20'h057ec: out <= 12'h000;
      20'h057ed: out <= 12'h000;
      20'h057ee: out <= 12'h000;
      20'h057ef: out <= 12'h000;
      20'h057f0: out <= 12'h222;
      20'h057f1: out <= 12'h222;
      20'h057f2: out <= 12'h222;
      20'h057f3: out <= 12'h222;
      20'h057f4: out <= 12'h222;
      20'h057f5: out <= 12'h222;
      20'h057f6: out <= 12'h222;
      20'h057f7: out <= 12'h222;
      20'h057f8: out <= 12'h222;
      20'h057f9: out <= 12'h222;
      20'h057fa: out <= 12'h222;
      20'h057fb: out <= 12'h222;
      20'h057fc: out <= 12'h222;
      20'h057fd: out <= 12'h222;
      20'h057fe: out <= 12'h222;
      20'h057ff: out <= 12'h222;
      20'h05800: out <= 12'h603;
      20'h05801: out <= 12'h603;
      20'h05802: out <= 12'h603;
      20'h05803: out <= 12'h603;
      20'h05804: out <= 12'hee9;
      20'h05805: out <= 12'hee9;
      20'h05806: out <= 12'hee9;
      20'h05807: out <= 12'hee9;
      20'h05808: out <= 12'hb27;
      20'h05809: out <= 12'hee9;
      20'h0580a: out <= 12'hee9;
      20'h0580b: out <= 12'hee9;
      20'h0580c: out <= 12'h000;
      20'h0580d: out <= 12'h000;
      20'h0580e: out <= 12'h000;
      20'h0580f: out <= 12'h000;
      20'h05810: out <= 12'hb27;
      20'h05811: out <= 12'hee9;
      20'h05812: out <= 12'hee9;
      20'h05813: out <= 12'hee9;
      20'h05814: out <= 12'h000;
      20'h05815: out <= 12'h000;
      20'h05816: out <= 12'h000;
      20'h05817: out <= 12'h000;
      20'h05818: out <= 12'h000;
      20'h05819: out <= 12'h000;
      20'h0581a: out <= 12'h000;
      20'h0581b: out <= 12'h000;
      20'h0581c: out <= 12'hee9;
      20'h0581d: out <= 12'hee9;
      20'h0581e: out <= 12'hee9;
      20'h0581f: out <= 12'hee9;
      20'h05820: out <= 12'h000;
      20'h05821: out <= 12'h000;
      20'h05822: out <= 12'h000;
      20'h05823: out <= 12'h000;
      20'h05824: out <= 12'hee9;
      20'h05825: out <= 12'hee9;
      20'h05826: out <= 12'hee9;
      20'h05827: out <= 12'hee9;
      20'h05828: out <= 12'hb27;
      20'h05829: out <= 12'hee9;
      20'h0582a: out <= 12'hee9;
      20'h0582b: out <= 12'hee9;
      20'h0582c: out <= 12'h603;
      20'h0582d: out <= 12'h603;
      20'h0582e: out <= 12'h603;
      20'h0582f: out <= 12'h603;
      20'h05830: out <= 12'h603;
      20'h05831: out <= 12'h603;
      20'h05832: out <= 12'h603;
      20'h05833: out <= 12'h603;
      20'h05834: out <= 12'hfff;
      20'h05835: out <= 12'hfff;
      20'h05836: out <= 12'hfff;
      20'h05837: out <= 12'hfff;
      20'h05838: out <= 12'hfff;
      20'h05839: out <= 12'hfff;
      20'h0583a: out <= 12'hfff;
      20'h0583b: out <= 12'h666;
      20'h0583c: out <= 12'h000;
      20'h0583d: out <= 12'h000;
      20'h0583e: out <= 12'hfff;
      20'h0583f: out <= 12'hfff;
      20'h05840: out <= 12'hfff;
      20'h05841: out <= 12'h8d0;
      20'h05842: out <= 12'h380;
      20'h05843: out <= 12'h000;
      20'h05844: out <= 12'hfff;
      20'h05845: out <= 12'h666;
      20'h05846: out <= 12'h000;
      20'h05847: out <= 12'h000;
      20'h05848: out <= 12'hfff;
      20'h05849: out <= 12'h666;
      20'h0584a: out <= 12'h000;
      20'h0584b: out <= 12'h000;
      20'h0584c: out <= 12'hfff;
      20'h0584d: out <= 12'h6af;
      20'h0584e: out <= 12'h6af;
      20'h0584f: out <= 12'hfff;
      20'h05850: out <= 12'h4cd;
      20'h05851: out <= 12'h4cd;
      20'h05852: out <= 12'h4cd;
      20'h05853: out <= 12'h4cd;
      20'h05854: out <= 12'h603;
      20'h05855: out <= 12'h603;
      20'h05856: out <= 12'h603;
      20'h05857: out <= 12'h603;
      20'h05858: out <= 12'hee9;
      20'h05859: out <= 12'hee9;
      20'h0585a: out <= 12'hee9;
      20'h0585b: out <= 12'hee9;
      20'h0585c: out <= 12'hee9;
      20'h0585d: out <= 12'hee9;
      20'h0585e: out <= 12'hee9;
      20'h0585f: out <= 12'hb27;
      20'h05860: out <= 12'h000;
      20'h05861: out <= 12'h000;
      20'h05862: out <= 12'h000;
      20'h05863: out <= 12'h000;
      20'h05864: out <= 12'h000;
      20'h05865: out <= 12'h000;
      20'h05866: out <= 12'h000;
      20'h05867: out <= 12'h000;
      20'h05868: out <= 12'h000;
      20'h05869: out <= 12'h6af;
      20'h0586a: out <= 12'hfff;
      20'h0586b: out <= 12'h16d;
      20'h0586c: out <= 12'h6af;
      20'h0586d: out <= 12'h16d;
      20'h0586e: out <= 12'h6af;
      20'h0586f: out <= 12'hfff;
      20'h05870: out <= 12'hfff;
      20'h05871: out <= 12'hfff;
      20'h05872: out <= 12'h6af;
      20'h05873: out <= 12'h16d;
      20'h05874: out <= 12'h6af;
      20'h05875: out <= 12'h16d;
      20'h05876: out <= 12'hfff;
      20'h05877: out <= 12'h6af;
      20'h05878: out <= 12'h000;
      20'h05879: out <= 12'h000;
      20'h0587a: out <= 12'h000;
      20'h0587b: out <= 12'h000;
      20'h0587c: out <= 12'h000;
      20'h0587d: out <= 12'h000;
      20'h0587e: out <= 12'h000;
      20'h0587f: out <= 12'h000;
      20'h05880: out <= 12'h4cd;
      20'h05881: out <= 12'h4cd;
      20'h05882: out <= 12'h4cd;
      20'h05883: out <= 12'h4cd;
      20'h05884: out <= 12'h4cd;
      20'h05885: out <= 12'h4cd;
      20'h05886: out <= 12'h4cd;
      20'h05887: out <= 12'h4cd;
      20'h05888: out <= 12'h5ef;
      20'h05889: out <= 12'h5ef;
      20'h0588a: out <= 12'h5ef;
      20'h0588b: out <= 12'h5ef;
      20'h0588c: out <= 12'h5ef;
      20'h0588d: out <= 12'h5ef;
      20'h0588e: out <= 12'h5ef;
      20'h0588f: out <= 12'h5ef;
      20'h05890: out <= 12'h000;
      20'h05891: out <= 12'h000;
      20'h05892: out <= 12'h000;
      20'h05893: out <= 12'h000;
      20'h05894: out <= 12'h000;
      20'h05895: out <= 12'h000;
      20'h05896: out <= 12'h000;
      20'h05897: out <= 12'h000;
      20'h05898: out <= 12'h000;
      20'h05899: out <= 12'h000;
      20'h0589a: out <= 12'h000;
      20'h0589b: out <= 12'h000;
      20'h0589c: out <= 12'h000;
      20'h0589d: out <= 12'h000;
      20'h0589e: out <= 12'h000;
      20'h0589f: out <= 12'h000;
      20'h058a0: out <= 12'h000;
      20'h058a1: out <= 12'h000;
      20'h058a2: out <= 12'h000;
      20'h058a3: out <= 12'h000;
      20'h058a4: out <= 12'h000;
      20'h058a5: out <= 12'h000;
      20'h058a6: out <= 12'h000;
      20'h058a7: out <= 12'h000;
      20'h058a8: out <= 12'h222;
      20'h058a9: out <= 12'h222;
      20'h058aa: out <= 12'h222;
      20'h058ab: out <= 12'h222;
      20'h058ac: out <= 12'h222;
      20'h058ad: out <= 12'h222;
      20'h058ae: out <= 12'h222;
      20'h058af: out <= 12'h222;
      20'h058b0: out <= 12'h222;
      20'h058b1: out <= 12'h222;
      20'h058b2: out <= 12'h222;
      20'h058b3: out <= 12'h222;
      20'h058b4: out <= 12'h222;
      20'h058b5: out <= 12'h222;
      20'h058b6: out <= 12'h222;
      20'h058b7: out <= 12'h222;
      20'h058b8: out <= 12'h000;
      20'h058b9: out <= 12'h000;
      20'h058ba: out <= 12'h000;
      20'h058bb: out <= 12'h000;
      20'h058bc: out <= 12'h000;
      20'h058bd: out <= 12'h000;
      20'h058be: out <= 12'h000;
      20'h058bf: out <= 12'h666;
      20'h058c0: out <= 12'hfff;
      20'h058c1: out <= 12'h666;
      20'h058c2: out <= 12'h000;
      20'h058c3: out <= 12'h000;
      20'h058c4: out <= 12'h000;
      20'h058c5: out <= 12'h000;
      20'h058c6: out <= 12'h000;
      20'h058c7: out <= 12'h000;
      20'h058c8: out <= 12'h222;
      20'h058c9: out <= 12'h222;
      20'h058ca: out <= 12'h222;
      20'h058cb: out <= 12'h222;
      20'h058cc: out <= 12'h222;
      20'h058cd: out <= 12'h222;
      20'h058ce: out <= 12'h222;
      20'h058cf: out <= 12'h666;
      20'h058d0: out <= 12'hfff;
      20'h058d1: out <= 12'h666;
      20'h058d2: out <= 12'h222;
      20'h058d3: out <= 12'h222;
      20'h058d4: out <= 12'h222;
      20'h058d5: out <= 12'h222;
      20'h058d6: out <= 12'h222;
      20'h058d7: out <= 12'h222;
      20'h058d8: out <= 12'h000;
      20'h058d9: out <= 12'h000;
      20'h058da: out <= 12'h000;
      20'h058db: out <= 12'h000;
      20'h058dc: out <= 12'h000;
      20'h058dd: out <= 12'h000;
      20'h058de: out <= 12'h000;
      20'h058df: out <= 12'h000;
      20'h058e0: out <= 12'h000;
      20'h058e1: out <= 12'h000;
      20'h058e2: out <= 12'h000;
      20'h058e3: out <= 12'h000;
      20'h058e4: out <= 12'h000;
      20'h058e5: out <= 12'h000;
      20'h058e6: out <= 12'h000;
      20'h058e7: out <= 12'h000;
      20'h058e8: out <= 12'h222;
      20'h058e9: out <= 12'h222;
      20'h058ea: out <= 12'h222;
      20'h058eb: out <= 12'h222;
      20'h058ec: out <= 12'h222;
      20'h058ed: out <= 12'h222;
      20'h058ee: out <= 12'h222;
      20'h058ef: out <= 12'h222;
      20'h058f0: out <= 12'h222;
      20'h058f1: out <= 12'h222;
      20'h058f2: out <= 12'h222;
      20'h058f3: out <= 12'h222;
      20'h058f4: out <= 12'h222;
      20'h058f5: out <= 12'h222;
      20'h058f6: out <= 12'h222;
      20'h058f7: out <= 12'h222;
      20'h058f8: out <= 12'h000;
      20'h058f9: out <= 12'h000;
      20'h058fa: out <= 12'h000;
      20'h058fb: out <= 12'h000;
      20'h058fc: out <= 12'h000;
      20'h058fd: out <= 12'h000;
      20'h058fe: out <= 12'h666;
      20'h058ff: out <= 12'h666;
      20'h05900: out <= 12'h666;
      20'h05901: out <= 12'h666;
      20'h05902: out <= 12'h666;
      20'h05903: out <= 12'h000;
      20'h05904: out <= 12'h000;
      20'h05905: out <= 12'h000;
      20'h05906: out <= 12'h000;
      20'h05907: out <= 12'h000;
      20'h05908: out <= 12'h222;
      20'h05909: out <= 12'h222;
      20'h0590a: out <= 12'h222;
      20'h0590b: out <= 12'h222;
      20'h0590c: out <= 12'h222;
      20'h0590d: out <= 12'h222;
      20'h0590e: out <= 12'h666;
      20'h0590f: out <= 12'h666;
      20'h05910: out <= 12'h666;
      20'h05911: out <= 12'h666;
      20'h05912: out <= 12'h666;
      20'h05913: out <= 12'h222;
      20'h05914: out <= 12'h222;
      20'h05915: out <= 12'h222;
      20'h05916: out <= 12'h222;
      20'h05917: out <= 12'h222;
      20'h05918: out <= 12'h603;
      20'h05919: out <= 12'h603;
      20'h0591a: out <= 12'h603;
      20'h0591b: out <= 12'h603;
      20'h0591c: out <= 12'hf87;
      20'h0591d: out <= 12'hf87;
      20'h0591e: out <= 12'hf87;
      20'h0591f: out <= 12'hee9;
      20'h05920: out <= 12'hb27;
      20'h05921: out <= 12'hf87;
      20'h05922: out <= 12'hf87;
      20'h05923: out <= 12'hf87;
      20'h05924: out <= 12'h000;
      20'h05925: out <= 12'h000;
      20'h05926: out <= 12'h000;
      20'h05927: out <= 12'h000;
      20'h05928: out <= 12'hb27;
      20'h05929: out <= 12'hf87;
      20'h0592a: out <= 12'hf87;
      20'h0592b: out <= 12'hf87;
      20'h0592c: out <= 12'h000;
      20'h0592d: out <= 12'h000;
      20'h0592e: out <= 12'h000;
      20'h0592f: out <= 12'h000;
      20'h05930: out <= 12'h000;
      20'h05931: out <= 12'h000;
      20'h05932: out <= 12'h000;
      20'h05933: out <= 12'h000;
      20'h05934: out <= 12'hf87;
      20'h05935: out <= 12'hf87;
      20'h05936: out <= 12'hf87;
      20'h05937: out <= 12'hee9;
      20'h05938: out <= 12'h000;
      20'h05939: out <= 12'h000;
      20'h0593a: out <= 12'h000;
      20'h0593b: out <= 12'h000;
      20'h0593c: out <= 12'hf87;
      20'h0593d: out <= 12'hf87;
      20'h0593e: out <= 12'hf87;
      20'h0593f: out <= 12'hee9;
      20'h05940: out <= 12'hb27;
      20'h05941: out <= 12'hf87;
      20'h05942: out <= 12'hf87;
      20'h05943: out <= 12'hf87;
      20'h05944: out <= 12'h603;
      20'h05945: out <= 12'h603;
      20'h05946: out <= 12'h603;
      20'h05947: out <= 12'h603;
      20'h05948: out <= 12'h603;
      20'h05949: out <= 12'h603;
      20'h0594a: out <= 12'h603;
      20'h0594b: out <= 12'h603;
      20'h0594c: out <= 12'hfff;
      20'h0594d: out <= 12'hbbb;
      20'h0594e: out <= 12'hbbb;
      20'h0594f: out <= 12'hbbb;
      20'h05950: out <= 12'hbbb;
      20'h05951: out <= 12'hbbb;
      20'h05952: out <= 12'h666;
      20'h05953: out <= 12'h666;
      20'h05954: out <= 12'h000;
      20'h05955: out <= 12'hfff;
      20'h05956: out <= 12'h8d0;
      20'h05957: out <= 12'hfff;
      20'h05958: out <= 12'h8d0;
      20'h05959: out <= 12'h380;
      20'h0595a: out <= 12'h8d0;
      20'h0595b: out <= 12'h380;
      20'h0595c: out <= 12'hbbb;
      20'h0595d: out <= 12'hfff;
      20'h0595e: out <= 12'h000;
      20'h0595f: out <= 12'h000;
      20'h05960: out <= 12'hbbb;
      20'h05961: out <= 12'hfff;
      20'h05962: out <= 12'h000;
      20'h05963: out <= 12'h000;
      20'h05964: out <= 12'h4cd;
      20'h05965: out <= 12'hfff;
      20'h05966: out <= 12'hfff;
      20'h05967: out <= 12'h4cd;
      20'h05968: out <= 12'h4cd;
      20'h05969: out <= 12'h6af;
      20'h0596a: out <= 12'h6af;
      20'h0596b: out <= 12'h4cd;
      20'h0596c: out <= 12'h603;
      20'h0596d: out <= 12'h603;
      20'h0596e: out <= 12'h603;
      20'h0596f: out <= 12'h603;
      20'h05970: out <= 12'hee9;
      20'h05971: out <= 12'hf87;
      20'h05972: out <= 12'hf87;
      20'h05973: out <= 12'hf87;
      20'h05974: out <= 12'hf87;
      20'h05975: out <= 12'hf87;
      20'h05976: out <= 12'hf87;
      20'h05977: out <= 12'hb27;
      20'h05978: out <= 12'h000;
      20'h05979: out <= 12'h000;
      20'h0597a: out <= 12'h000;
      20'h0597b: out <= 12'h000;
      20'h0597c: out <= 12'h000;
      20'h0597d: out <= 12'h000;
      20'h0597e: out <= 12'h000;
      20'h0597f: out <= 12'h000;
      20'h05980: out <= 12'h000;
      20'h05981: out <= 12'h6af;
      20'h05982: out <= 12'h16d;
      20'h05983: out <= 12'h16d;
      20'h05984: out <= 12'h6af;
      20'h05985: out <= 12'h16d;
      20'h05986: out <= 12'h16d;
      20'h05987: out <= 12'h6af;
      20'h05988: out <= 12'hfff;
      20'h05989: out <= 12'h6af;
      20'h0598a: out <= 12'h16d;
      20'h0598b: out <= 12'h16d;
      20'h0598c: out <= 12'h6af;
      20'h0598d: out <= 12'h16d;
      20'h0598e: out <= 12'h16d;
      20'h0598f: out <= 12'h6af;
      20'h05990: out <= 12'h000;
      20'h05991: out <= 12'h000;
      20'h05992: out <= 12'h4cd;
      20'h05993: out <= 12'h000;
      20'h05994: out <= 12'h000;
      20'h05995: out <= 12'h000;
      20'h05996: out <= 12'h4cd;
      20'h05997: out <= 12'h000;
      20'h05998: out <= 12'h4cd;
      20'h05999: out <= 12'h4cd;
      20'h0599a: out <= 12'h4cd;
      20'h0599b: out <= 12'h4cd;
      20'h0599c: out <= 12'h4cd;
      20'h0599d: out <= 12'h4cd;
      20'h0599e: out <= 12'h4cd;
      20'h0599f: out <= 12'h4cd;
      20'h059a0: out <= 12'h5ef;
      20'h059a1: out <= 12'h5ef;
      20'h059a2: out <= 12'h5ef;
      20'h059a3: out <= 12'h5ef;
      20'h059a4: out <= 12'h5ef;
      20'h059a5: out <= 12'h5ef;
      20'h059a6: out <= 12'h5ef;
      20'h059a7: out <= 12'h5ef;
      20'h059a8: out <= 12'h000;
      20'h059a9: out <= 12'h000;
      20'h059aa: out <= 12'h000;
      20'h059ab: out <= 12'h000;
      20'h059ac: out <= 12'h000;
      20'h059ad: out <= 12'h000;
      20'h059ae: out <= 12'h000;
      20'h059af: out <= 12'h000;
      20'h059b0: out <= 12'h000;
      20'h059b1: out <= 12'h000;
      20'h059b2: out <= 12'h000;
      20'h059b3: out <= 12'hfff;
      20'h059b4: out <= 12'h666;
      20'h059b5: out <= 12'hbbb;
      20'h059b6: out <= 12'h666;
      20'h059b7: out <= 12'hbbb;
      20'h059b8: out <= 12'h666;
      20'h059b9: out <= 12'hbbb;
      20'h059ba: out <= 12'h666;
      20'h059bb: out <= 12'hfff;
      20'h059bc: out <= 12'h000;
      20'h059bd: out <= 12'h000;
      20'h059be: out <= 12'h000;
      20'h059bf: out <= 12'h000;
      20'h059c0: out <= 12'h222;
      20'h059c1: out <= 12'h222;
      20'h059c2: out <= 12'h222;
      20'h059c3: out <= 12'hfff;
      20'h059c4: out <= 12'hbbb;
      20'h059c5: out <= 12'h666;
      20'h059c6: out <= 12'hbbb;
      20'h059c7: out <= 12'h666;
      20'h059c8: out <= 12'hbbb;
      20'h059c9: out <= 12'h666;
      20'h059ca: out <= 12'hbbb;
      20'h059cb: out <= 12'hfff;
      20'h059cc: out <= 12'h222;
      20'h059cd: out <= 12'h222;
      20'h059ce: out <= 12'h222;
      20'h059cf: out <= 12'h222;
      20'h059d0: out <= 12'h000;
      20'h059d1: out <= 12'h000;
      20'h059d2: out <= 12'h000;
      20'h059d3: out <= 12'h000;
      20'h059d4: out <= 12'h000;
      20'h059d5: out <= 12'h000;
      20'h059d6: out <= 12'h000;
      20'h059d7: out <= 12'h666;
      20'h059d8: out <= 12'hfff;
      20'h059d9: out <= 12'h666;
      20'h059da: out <= 12'h000;
      20'h059db: out <= 12'h000;
      20'h059dc: out <= 12'h000;
      20'h059dd: out <= 12'h000;
      20'h059de: out <= 12'h000;
      20'h059df: out <= 12'h000;
      20'h059e0: out <= 12'h222;
      20'h059e1: out <= 12'h222;
      20'h059e2: out <= 12'h222;
      20'h059e3: out <= 12'h222;
      20'h059e4: out <= 12'h222;
      20'h059e5: out <= 12'h222;
      20'h059e6: out <= 12'h222;
      20'h059e7: out <= 12'h666;
      20'h059e8: out <= 12'hfff;
      20'h059e9: out <= 12'h666;
      20'h059ea: out <= 12'h222;
      20'h059eb: out <= 12'h222;
      20'h059ec: out <= 12'h222;
      20'h059ed: out <= 12'h222;
      20'h059ee: out <= 12'h222;
      20'h059ef: out <= 12'h222;
      20'h059f0: out <= 12'h000;
      20'h059f1: out <= 12'h000;
      20'h059f2: out <= 12'h000;
      20'h059f3: out <= 12'h000;
      20'h059f4: out <= 12'hfff;
      20'h059f5: out <= 12'h666;
      20'h059f6: out <= 12'hbbb;
      20'h059f7: out <= 12'h666;
      20'h059f8: out <= 12'hbbb;
      20'h059f9: out <= 12'h666;
      20'h059fa: out <= 12'hbbb;
      20'h059fb: out <= 12'h666;
      20'h059fc: out <= 12'hfff;
      20'h059fd: out <= 12'h000;
      20'h059fe: out <= 12'h000;
      20'h059ff: out <= 12'h000;
      20'h05a00: out <= 12'h222;
      20'h05a01: out <= 12'h222;
      20'h05a02: out <= 12'h222;
      20'h05a03: out <= 12'h222;
      20'h05a04: out <= 12'hfff;
      20'h05a05: out <= 12'hbbb;
      20'h05a06: out <= 12'h666;
      20'h05a07: out <= 12'hbbb;
      20'h05a08: out <= 12'h666;
      20'h05a09: out <= 12'hbbb;
      20'h05a0a: out <= 12'h666;
      20'h05a0b: out <= 12'hbbb;
      20'h05a0c: out <= 12'hfff;
      20'h05a0d: out <= 12'h222;
      20'h05a0e: out <= 12'h222;
      20'h05a0f: out <= 12'h222;
      20'h05a10: out <= 12'h000;
      20'h05a11: out <= 12'h000;
      20'h05a12: out <= 12'h000;
      20'h05a13: out <= 12'h000;
      20'h05a14: out <= 12'h000;
      20'h05a15: out <= 12'h666;
      20'h05a16: out <= 12'hbbb;
      20'h05a17: out <= 12'hbbb;
      20'h05a18: out <= 12'hbbb;
      20'h05a19: out <= 12'hbbb;
      20'h05a1a: out <= 12'hbbb;
      20'h05a1b: out <= 12'h666;
      20'h05a1c: out <= 12'h000;
      20'h05a1d: out <= 12'h000;
      20'h05a1e: out <= 12'h000;
      20'h05a1f: out <= 12'h000;
      20'h05a20: out <= 12'h222;
      20'h05a21: out <= 12'h222;
      20'h05a22: out <= 12'h222;
      20'h05a23: out <= 12'h222;
      20'h05a24: out <= 12'h222;
      20'h05a25: out <= 12'h666;
      20'h05a26: out <= 12'hbbb;
      20'h05a27: out <= 12'hbbb;
      20'h05a28: out <= 12'hbbb;
      20'h05a29: out <= 12'hbbb;
      20'h05a2a: out <= 12'hbbb;
      20'h05a2b: out <= 12'h666;
      20'h05a2c: out <= 12'h222;
      20'h05a2d: out <= 12'h222;
      20'h05a2e: out <= 12'h222;
      20'h05a2f: out <= 12'h222;
      20'h05a30: out <= 12'h603;
      20'h05a31: out <= 12'h603;
      20'h05a32: out <= 12'h603;
      20'h05a33: out <= 12'h603;
      20'h05a34: out <= 12'hf87;
      20'h05a35: out <= 12'hf87;
      20'h05a36: out <= 12'hf87;
      20'h05a37: out <= 12'hee9;
      20'h05a38: out <= 12'hb27;
      20'h05a39: out <= 12'hf87;
      20'h05a3a: out <= 12'hf87;
      20'h05a3b: out <= 12'hf87;
      20'h05a3c: out <= 12'h000;
      20'h05a3d: out <= 12'h000;
      20'h05a3e: out <= 12'h000;
      20'h05a3f: out <= 12'h000;
      20'h05a40: out <= 12'hb27;
      20'h05a41: out <= 12'hf87;
      20'h05a42: out <= 12'hf87;
      20'h05a43: out <= 12'hf87;
      20'h05a44: out <= 12'h000;
      20'h05a45: out <= 12'h000;
      20'h05a46: out <= 12'h000;
      20'h05a47: out <= 12'h000;
      20'h05a48: out <= 12'h000;
      20'h05a49: out <= 12'h000;
      20'h05a4a: out <= 12'h000;
      20'h05a4b: out <= 12'h000;
      20'h05a4c: out <= 12'hf87;
      20'h05a4d: out <= 12'hf87;
      20'h05a4e: out <= 12'hf87;
      20'h05a4f: out <= 12'hee9;
      20'h05a50: out <= 12'h000;
      20'h05a51: out <= 12'h000;
      20'h05a52: out <= 12'h000;
      20'h05a53: out <= 12'h000;
      20'h05a54: out <= 12'hf87;
      20'h05a55: out <= 12'hf87;
      20'h05a56: out <= 12'hf87;
      20'h05a57: out <= 12'hee9;
      20'h05a58: out <= 12'hb27;
      20'h05a59: out <= 12'hf87;
      20'h05a5a: out <= 12'hf87;
      20'h05a5b: out <= 12'hf87;
      20'h05a5c: out <= 12'h603;
      20'h05a5d: out <= 12'h603;
      20'h05a5e: out <= 12'h603;
      20'h05a5f: out <= 12'h603;
      20'h05a60: out <= 12'h603;
      20'h05a61: out <= 12'h603;
      20'h05a62: out <= 12'h603;
      20'h05a63: out <= 12'h603;
      20'h05a64: out <= 12'hfff;
      20'h05a65: out <= 12'hbbb;
      20'h05a66: out <= 12'h666;
      20'h05a67: out <= 12'h666;
      20'h05a68: out <= 12'h666;
      20'h05a69: out <= 12'hbbb;
      20'h05a6a: out <= 12'h666;
      20'h05a6b: out <= 12'h666;
      20'h05a6c: out <= 12'hfff;
      20'h05a6d: out <= 12'h8d0;
      20'h05a6e: out <= 12'hfff;
      20'h05a6f: out <= 12'h8d0;
      20'h05a70: out <= 12'h8d0;
      20'h05a71: out <= 12'h8d0;
      20'h05a72: out <= 12'h380;
      20'h05a73: out <= 12'h8d0;
      20'h05a74: out <= 12'h000;
      20'h05a75: out <= 12'h000;
      20'h05a76: out <= 12'hfff;
      20'h05a77: out <= 12'h666;
      20'h05a78: out <= 12'h000;
      20'h05a79: out <= 12'h000;
      20'h05a7a: out <= 12'hfff;
      20'h05a7b: out <= 12'h666;
      20'h05a7c: out <= 12'h4cd;
      20'h05a7d: out <= 12'h4cd;
      20'h05a7e: out <= 12'h4cd;
      20'h05a7f: out <= 12'h4cd;
      20'h05a80: out <= 12'h6af;
      20'h05a81: out <= 12'hfff;
      20'h05a82: out <= 12'hfff;
      20'h05a83: out <= 12'h6af;
      20'h05a84: out <= 12'h603;
      20'h05a85: out <= 12'h603;
      20'h05a86: out <= 12'h603;
      20'h05a87: out <= 12'h603;
      20'h05a88: out <= 12'hee9;
      20'h05a89: out <= 12'hf87;
      20'h05a8a: out <= 12'hee9;
      20'h05a8b: out <= 12'hee9;
      20'h05a8c: out <= 12'hee9;
      20'h05a8d: out <= 12'hb27;
      20'h05a8e: out <= 12'hf87;
      20'h05a8f: out <= 12'hb27;
      20'h05a90: out <= 12'h000;
      20'h05a91: out <= 12'h000;
      20'h05a92: out <= 12'h000;
      20'h05a93: out <= 12'h000;
      20'h05a94: out <= 12'h000;
      20'h05a95: out <= 12'h000;
      20'h05a96: out <= 12'h000;
      20'h05a97: out <= 12'h000;
      20'h05a98: out <= 12'h000;
      20'h05a99: out <= 12'h6af;
      20'h05a9a: out <= 12'hfff;
      20'h05a9b: out <= 12'h16d;
      20'h05a9c: out <= 12'h6af;
      20'h05a9d: out <= 12'h6af;
      20'h05a9e: out <= 12'h16d;
      20'h05a9f: out <= 12'h16d;
      20'h05aa0: out <= 12'h6af;
      20'h05aa1: out <= 12'h16d;
      20'h05aa2: out <= 12'h16d;
      20'h05aa3: out <= 12'h6af;
      20'h05aa4: out <= 12'h6af;
      20'h05aa5: out <= 12'h16d;
      20'h05aa6: out <= 12'hfff;
      20'h05aa7: out <= 12'h6af;
      20'h05aa8: out <= 12'h000;
      20'h05aa9: out <= 12'h000;
      20'h05aaa: out <= 12'h000;
      20'h05aab: out <= 12'h4cd;
      20'h05aac: out <= 12'h000;
      20'h05aad: out <= 12'h4cd;
      20'h05aae: out <= 12'h000;
      20'h05aaf: out <= 12'h000;
      20'h05ab0: out <= 12'h4cd;
      20'h05ab1: out <= 12'h4cd;
      20'h05ab2: out <= 12'h4cd;
      20'h05ab3: out <= 12'h4cd;
      20'h05ab4: out <= 12'h4cd;
      20'h05ab5: out <= 12'h4cd;
      20'h05ab6: out <= 12'h4cd;
      20'h05ab7: out <= 12'h4cd;
      20'h05ab8: out <= 12'h5ef;
      20'h05ab9: out <= 12'h5ef;
      20'h05aba: out <= 12'h5ef;
      20'h05abb: out <= 12'h5ef;
      20'h05abc: out <= 12'h5ef;
      20'h05abd: out <= 12'h5ef;
      20'h05abe: out <= 12'h5ef;
      20'h05abf: out <= 12'h5ef;
      20'h05ac0: out <= 12'h000;
      20'h05ac1: out <= 12'h000;
      20'h05ac2: out <= 12'h000;
      20'h05ac3: out <= 12'h000;
      20'h05ac4: out <= 12'h000;
      20'h05ac5: out <= 12'h000;
      20'h05ac6: out <= 12'h000;
      20'h05ac7: out <= 12'h000;
      20'h05ac8: out <= 12'h000;
      20'h05ac9: out <= 12'h000;
      20'h05aca: out <= 12'h000;
      20'h05acb: out <= 12'h666;
      20'h05acc: out <= 12'h666;
      20'h05acd: out <= 12'h666;
      20'h05ace: out <= 12'h666;
      20'h05acf: out <= 12'h666;
      20'h05ad0: out <= 12'h666;
      20'h05ad1: out <= 12'h666;
      20'h05ad2: out <= 12'h666;
      20'h05ad3: out <= 12'h666;
      20'h05ad4: out <= 12'h000;
      20'h05ad5: out <= 12'h000;
      20'h05ad6: out <= 12'h000;
      20'h05ad7: out <= 12'h000;
      20'h05ad8: out <= 12'h222;
      20'h05ad9: out <= 12'h222;
      20'h05ada: out <= 12'h222;
      20'h05adb: out <= 12'h666;
      20'h05adc: out <= 12'h666;
      20'h05add: out <= 12'h666;
      20'h05ade: out <= 12'h666;
      20'h05adf: out <= 12'h666;
      20'h05ae0: out <= 12'h666;
      20'h05ae1: out <= 12'h666;
      20'h05ae2: out <= 12'h666;
      20'h05ae3: out <= 12'h666;
      20'h05ae4: out <= 12'h222;
      20'h05ae5: out <= 12'h222;
      20'h05ae6: out <= 12'h222;
      20'h05ae7: out <= 12'h222;
      20'h05ae8: out <= 12'h000;
      20'h05ae9: out <= 12'h000;
      20'h05aea: out <= 12'h000;
      20'h05aeb: out <= 12'h000;
      20'h05aec: out <= 12'h000;
      20'h05aed: out <= 12'h666;
      20'h05aee: out <= 12'h666;
      20'h05aef: out <= 12'h666;
      20'h05af0: out <= 12'hfff;
      20'h05af1: out <= 12'h666;
      20'h05af2: out <= 12'h666;
      20'h05af3: out <= 12'h666;
      20'h05af4: out <= 12'h000;
      20'h05af5: out <= 12'h000;
      20'h05af6: out <= 12'h000;
      20'h05af7: out <= 12'h000;
      20'h05af8: out <= 12'h222;
      20'h05af9: out <= 12'h222;
      20'h05afa: out <= 12'h222;
      20'h05afb: out <= 12'h222;
      20'h05afc: out <= 12'h222;
      20'h05afd: out <= 12'h666;
      20'h05afe: out <= 12'h666;
      20'h05aff: out <= 12'h666;
      20'h05b00: out <= 12'hfff;
      20'h05b01: out <= 12'h666;
      20'h05b02: out <= 12'h666;
      20'h05b03: out <= 12'h666;
      20'h05b04: out <= 12'h222;
      20'h05b05: out <= 12'h222;
      20'h05b06: out <= 12'h222;
      20'h05b07: out <= 12'h222;
      20'h05b08: out <= 12'h000;
      20'h05b09: out <= 12'h000;
      20'h05b0a: out <= 12'h000;
      20'h05b0b: out <= 12'h000;
      20'h05b0c: out <= 12'h666;
      20'h05b0d: out <= 12'h666;
      20'h05b0e: out <= 12'h666;
      20'h05b0f: out <= 12'h666;
      20'h05b10: out <= 12'h666;
      20'h05b11: out <= 12'h666;
      20'h05b12: out <= 12'h666;
      20'h05b13: out <= 12'h666;
      20'h05b14: out <= 12'h666;
      20'h05b15: out <= 12'h000;
      20'h05b16: out <= 12'h000;
      20'h05b17: out <= 12'h000;
      20'h05b18: out <= 12'h222;
      20'h05b19: out <= 12'h222;
      20'h05b1a: out <= 12'h222;
      20'h05b1b: out <= 12'h222;
      20'h05b1c: out <= 12'h666;
      20'h05b1d: out <= 12'h666;
      20'h05b1e: out <= 12'h666;
      20'h05b1f: out <= 12'h666;
      20'h05b20: out <= 12'h666;
      20'h05b21: out <= 12'h666;
      20'h05b22: out <= 12'h666;
      20'h05b23: out <= 12'h666;
      20'h05b24: out <= 12'h666;
      20'h05b25: out <= 12'h222;
      20'h05b26: out <= 12'h222;
      20'h05b27: out <= 12'h222;
      20'h05b28: out <= 12'h000;
      20'h05b29: out <= 12'h000;
      20'h05b2a: out <= 12'h000;
      20'h05b2b: out <= 12'hfff;
      20'h05b2c: out <= 12'h666;
      20'h05b2d: out <= 12'hbbb;
      20'h05b2e: out <= 12'hfff;
      20'h05b2f: out <= 12'h666;
      20'h05b30: out <= 12'h666;
      20'h05b31: out <= 12'h666;
      20'h05b32: out <= 12'h666;
      20'h05b33: out <= 12'hbbb;
      20'h05b34: out <= 12'h666;
      20'h05b35: out <= 12'hfff;
      20'h05b36: out <= 12'h000;
      20'h05b37: out <= 12'h000;
      20'h05b38: out <= 12'h222;
      20'h05b39: out <= 12'h222;
      20'h05b3a: out <= 12'h222;
      20'h05b3b: out <= 12'hfff;
      20'h05b3c: out <= 12'h666;
      20'h05b3d: out <= 12'hbbb;
      20'h05b3e: out <= 12'hfff;
      20'h05b3f: out <= 12'h666;
      20'h05b40: out <= 12'h666;
      20'h05b41: out <= 12'h666;
      20'h05b42: out <= 12'h666;
      20'h05b43: out <= 12'hbbb;
      20'h05b44: out <= 12'h666;
      20'h05b45: out <= 12'hfff;
      20'h05b46: out <= 12'h222;
      20'h05b47: out <= 12'h222;
      20'h05b48: out <= 12'h603;
      20'h05b49: out <= 12'h603;
      20'h05b4a: out <= 12'h603;
      20'h05b4b: out <= 12'h603;
      20'h05b4c: out <= 12'hb27;
      20'h05b4d: out <= 12'hb27;
      20'h05b4e: out <= 12'hb27;
      20'h05b4f: out <= 12'hb27;
      20'h05b50: out <= 12'hb27;
      20'h05b51: out <= 12'hb27;
      20'h05b52: out <= 12'hb27;
      20'h05b53: out <= 12'hb27;
      20'h05b54: out <= 12'h000;
      20'h05b55: out <= 12'h000;
      20'h05b56: out <= 12'h000;
      20'h05b57: out <= 12'h000;
      20'h05b58: out <= 12'hb27;
      20'h05b59: out <= 12'hb27;
      20'h05b5a: out <= 12'hb27;
      20'h05b5b: out <= 12'hb27;
      20'h05b5c: out <= 12'h000;
      20'h05b5d: out <= 12'h000;
      20'h05b5e: out <= 12'h000;
      20'h05b5f: out <= 12'h000;
      20'h05b60: out <= 12'h000;
      20'h05b61: out <= 12'h000;
      20'h05b62: out <= 12'h000;
      20'h05b63: out <= 12'h000;
      20'h05b64: out <= 12'hb27;
      20'h05b65: out <= 12'hb27;
      20'h05b66: out <= 12'hb27;
      20'h05b67: out <= 12'hb27;
      20'h05b68: out <= 12'h000;
      20'h05b69: out <= 12'h000;
      20'h05b6a: out <= 12'h000;
      20'h05b6b: out <= 12'h000;
      20'h05b6c: out <= 12'hb27;
      20'h05b6d: out <= 12'hb27;
      20'h05b6e: out <= 12'hb27;
      20'h05b6f: out <= 12'hb27;
      20'h05b70: out <= 12'hb27;
      20'h05b71: out <= 12'hb27;
      20'h05b72: out <= 12'hb27;
      20'h05b73: out <= 12'hb27;
      20'h05b74: out <= 12'h603;
      20'h05b75: out <= 12'h603;
      20'h05b76: out <= 12'h603;
      20'h05b77: out <= 12'h603;
      20'h05b78: out <= 12'h603;
      20'h05b79: out <= 12'h603;
      20'h05b7a: out <= 12'h603;
      20'h05b7b: out <= 12'h603;
      20'h05b7c: out <= 12'hfff;
      20'h05b7d: out <= 12'hbbb;
      20'h05b7e: out <= 12'h666;
      20'h05b7f: out <= 12'hbbb;
      20'h05b80: out <= 12'hfff;
      20'h05b81: out <= 12'hbbb;
      20'h05b82: out <= 12'h666;
      20'h05b83: out <= 12'h666;
      20'h05b84: out <= 12'h380;
      20'h05b85: out <= 12'hfff;
      20'h05b86: out <= 12'h8d0;
      20'h05b87: out <= 12'h8d0;
      20'h05b88: out <= 12'h380;
      20'h05b89: out <= 12'h000;
      20'h05b8a: out <= 12'h8d0;
      20'h05b8b: out <= 12'h000;
      20'h05b8c: out <= 12'h000;
      20'h05b8d: out <= 12'h000;
      20'h05b8e: out <= 12'hbbb;
      20'h05b8f: out <= 12'hfff;
      20'h05b90: out <= 12'h000;
      20'h05b91: out <= 12'h000;
      20'h05b92: out <= 12'hbbb;
      20'h05b93: out <= 12'hfff;
      20'h05b94: out <= 12'h6af;
      20'h05b95: out <= 12'h4cd;
      20'h05b96: out <= 12'h4cd;
      20'h05b97: out <= 12'h6af;
      20'h05b98: out <= 12'hfff;
      20'h05b99: out <= 12'h4cd;
      20'h05b9a: out <= 12'h4cd;
      20'h05b9b: out <= 12'hfff;
      20'h05b9c: out <= 12'h603;
      20'h05b9d: out <= 12'h603;
      20'h05b9e: out <= 12'h603;
      20'h05b9f: out <= 12'h603;
      20'h05ba0: out <= 12'hee9;
      20'h05ba1: out <= 12'hf87;
      20'h05ba2: out <= 12'hee9;
      20'h05ba3: out <= 12'hf87;
      20'h05ba4: out <= 12'hf87;
      20'h05ba5: out <= 12'hb27;
      20'h05ba6: out <= 12'hf87;
      20'h05ba7: out <= 12'hb27;
      20'h05ba8: out <= 12'h000;
      20'h05ba9: out <= 12'h000;
      20'h05baa: out <= 12'h000;
      20'h05bab: out <= 12'h000;
      20'h05bac: out <= 12'h000;
      20'h05bad: out <= 12'h000;
      20'h05bae: out <= 12'h000;
      20'h05baf: out <= 12'h000;
      20'h05bb0: out <= 12'h000;
      20'h05bb1: out <= 12'h6af;
      20'h05bb2: out <= 12'h16d;
      20'h05bb3: out <= 12'h16d;
      20'h05bb4: out <= 12'hfff;
      20'h05bb5: out <= 12'h6af;
      20'h05bb6: out <= 12'h6af;
      20'h05bb7: out <= 12'h16d;
      20'h05bb8: out <= 12'h16d;
      20'h05bb9: out <= 12'h16d;
      20'h05bba: out <= 12'h6af;
      20'h05bbb: out <= 12'h6af;
      20'h05bbc: out <= 12'hfff;
      20'h05bbd: out <= 12'h16d;
      20'h05bbe: out <= 12'h16d;
      20'h05bbf: out <= 12'h6af;
      20'h05bc0: out <= 12'h000;
      20'h05bc1: out <= 12'h000;
      20'h05bc2: out <= 12'h000;
      20'h05bc3: out <= 12'h000;
      20'h05bc4: out <= 12'h4cd;
      20'h05bc5: out <= 12'h000;
      20'h05bc6: out <= 12'h000;
      20'h05bc7: out <= 12'h000;
      20'h05bc8: out <= 12'h4cd;
      20'h05bc9: out <= 12'h4cd;
      20'h05bca: out <= 12'h4cd;
      20'h05bcb: out <= 12'h4cd;
      20'h05bcc: out <= 12'h4cd;
      20'h05bcd: out <= 12'h4cd;
      20'h05bce: out <= 12'h4cd;
      20'h05bcf: out <= 12'h4cd;
      20'h05bd0: out <= 12'h5ef;
      20'h05bd1: out <= 12'h5ef;
      20'h05bd2: out <= 12'h5ef;
      20'h05bd3: out <= 12'h5ef;
      20'h05bd4: out <= 12'h5ef;
      20'h05bd5: out <= 12'h5ef;
      20'h05bd6: out <= 12'h5ef;
      20'h05bd7: out <= 12'h5ef;
      20'h05bd8: out <= 12'h000;
      20'h05bd9: out <= 12'h000;
      20'h05bda: out <= 12'h000;
      20'h05bdb: out <= 12'h000;
      20'h05bdc: out <= 12'h000;
      20'h05bdd: out <= 12'h000;
      20'h05bde: out <= 12'h000;
      20'h05bdf: out <= 12'h000;
      20'h05be0: out <= 12'h000;
      20'h05be1: out <= 12'h000;
      20'h05be2: out <= 12'h666;
      20'h05be3: out <= 12'hbbb;
      20'h05be4: out <= 12'hbbb;
      20'h05be5: out <= 12'hbbb;
      20'h05be6: out <= 12'hbbb;
      20'h05be7: out <= 12'hbbb;
      20'h05be8: out <= 12'hbbb;
      20'h05be9: out <= 12'h666;
      20'h05bea: out <= 12'hbbb;
      20'h05beb: out <= 12'hfff;
      20'h05bec: out <= 12'h666;
      20'h05bed: out <= 12'h000;
      20'h05bee: out <= 12'h000;
      20'h05bef: out <= 12'h000;
      20'h05bf0: out <= 12'h222;
      20'h05bf1: out <= 12'h222;
      20'h05bf2: out <= 12'h666;
      20'h05bf3: out <= 12'hbbb;
      20'h05bf4: out <= 12'hbbb;
      20'h05bf5: out <= 12'hbbb;
      20'h05bf6: out <= 12'hbbb;
      20'h05bf7: out <= 12'hbbb;
      20'h05bf8: out <= 12'hbbb;
      20'h05bf9: out <= 12'h666;
      20'h05bfa: out <= 12'hbbb;
      20'h05bfb: out <= 12'hfff;
      20'h05bfc: out <= 12'h666;
      20'h05bfd: out <= 12'h222;
      20'h05bfe: out <= 12'h222;
      20'h05bff: out <= 12'h222;
      20'h05c00: out <= 12'h000;
      20'h05c01: out <= 12'h000;
      20'h05c02: out <= 12'h000;
      20'h05c03: out <= 12'hfff;
      20'h05c04: out <= 12'h666;
      20'h05c05: out <= 12'hfff;
      20'h05c06: out <= 12'hbbb;
      20'h05c07: out <= 12'h666;
      20'h05c08: out <= 12'hbbb;
      20'h05c09: out <= 12'h666;
      20'h05c0a: out <= 12'hbbb;
      20'h05c0b: out <= 12'hfff;
      20'h05c0c: out <= 12'h666;
      20'h05c0d: out <= 12'hfff;
      20'h05c0e: out <= 12'h000;
      20'h05c0f: out <= 12'h000;
      20'h05c10: out <= 12'h222;
      20'h05c11: out <= 12'h222;
      20'h05c12: out <= 12'h222;
      20'h05c13: out <= 12'hfff;
      20'h05c14: out <= 12'h666;
      20'h05c15: out <= 12'hfff;
      20'h05c16: out <= 12'hbbb;
      20'h05c17: out <= 12'h666;
      20'h05c18: out <= 12'hbbb;
      20'h05c19: out <= 12'h666;
      20'h05c1a: out <= 12'hbbb;
      20'h05c1b: out <= 12'hfff;
      20'h05c1c: out <= 12'h666;
      20'h05c1d: out <= 12'hfff;
      20'h05c1e: out <= 12'h222;
      20'h05c1f: out <= 12'h222;
      20'h05c20: out <= 12'h000;
      20'h05c21: out <= 12'h000;
      20'h05c22: out <= 12'h000;
      20'h05c23: out <= 12'h666;
      20'h05c24: out <= 12'hfff;
      20'h05c25: out <= 12'hbbb;
      20'h05c26: out <= 12'h666;
      20'h05c27: out <= 12'hbbb;
      20'h05c28: out <= 12'hbbb;
      20'h05c29: out <= 12'hbbb;
      20'h05c2a: out <= 12'hbbb;
      20'h05c2b: out <= 12'hbbb;
      20'h05c2c: out <= 12'hbbb;
      20'h05c2d: out <= 12'h666;
      20'h05c2e: out <= 12'h000;
      20'h05c2f: out <= 12'h000;
      20'h05c30: out <= 12'h222;
      20'h05c31: out <= 12'h222;
      20'h05c32: out <= 12'h222;
      20'h05c33: out <= 12'h666;
      20'h05c34: out <= 12'hfff;
      20'h05c35: out <= 12'hbbb;
      20'h05c36: out <= 12'h666;
      20'h05c37: out <= 12'hbbb;
      20'h05c38: out <= 12'hbbb;
      20'h05c39: out <= 12'hbbb;
      20'h05c3a: out <= 12'hbbb;
      20'h05c3b: out <= 12'hbbb;
      20'h05c3c: out <= 12'hbbb;
      20'h05c3d: out <= 12'h666;
      20'h05c3e: out <= 12'h222;
      20'h05c3f: out <= 12'h222;
      20'h05c40: out <= 12'h000;
      20'h05c41: out <= 12'h000;
      20'h05c42: out <= 12'h000;
      20'h05c43: out <= 12'h666;
      20'h05c44: out <= 12'h666;
      20'h05c45: out <= 12'hbbb;
      20'h05c46: out <= 12'hfff;
      20'h05c47: out <= 12'hbbb;
      20'h05c48: out <= 12'hbbb;
      20'h05c49: out <= 12'hbbb;
      20'h05c4a: out <= 12'h666;
      20'h05c4b: out <= 12'hbbb;
      20'h05c4c: out <= 12'h666;
      20'h05c4d: out <= 12'hbbb;
      20'h05c4e: out <= 12'h000;
      20'h05c4f: out <= 12'h000;
      20'h05c50: out <= 12'h222;
      20'h05c51: out <= 12'h222;
      20'h05c52: out <= 12'h222;
      20'h05c53: out <= 12'hbbb;
      20'h05c54: out <= 12'h666;
      20'h05c55: out <= 12'hbbb;
      20'h05c56: out <= 12'hfff;
      20'h05c57: out <= 12'hbbb;
      20'h05c58: out <= 12'hbbb;
      20'h05c59: out <= 12'hbbb;
      20'h05c5a: out <= 12'h666;
      20'h05c5b: out <= 12'hbbb;
      20'h05c5c: out <= 12'h666;
      20'h05c5d: out <= 12'h666;
      20'h05c5e: out <= 12'h222;
      20'h05c5f: out <= 12'h222;
      20'h05c60: out <= 12'h603;
      20'h05c61: out <= 12'h603;
      20'h05c62: out <= 12'h603;
      20'h05c63: out <= 12'h603;
      20'h05c64: out <= 12'hb27;
      20'h05c65: out <= 12'hee9;
      20'h05c66: out <= 12'hee9;
      20'h05c67: out <= 12'hee9;
      20'h05c68: out <= 12'hee9;
      20'h05c69: out <= 12'hee9;
      20'h05c6a: out <= 12'hee9;
      20'h05c6b: out <= 12'hee9;
      20'h05c6c: out <= 12'h000;
      20'h05c6d: out <= 12'h000;
      20'h05c6e: out <= 12'h000;
      20'h05c6f: out <= 12'h000;
      20'h05c70: out <= 12'hee9;
      20'h05c71: out <= 12'hee9;
      20'h05c72: out <= 12'hee9;
      20'h05c73: out <= 12'hee9;
      20'h05c74: out <= 12'hb27;
      20'h05c75: out <= 12'hee9;
      20'h05c76: out <= 12'hee9;
      20'h05c77: out <= 12'hee9;
      20'h05c78: out <= 12'hee9;
      20'h05c79: out <= 12'hee9;
      20'h05c7a: out <= 12'hee9;
      20'h05c7b: out <= 12'hee9;
      20'h05c7c: out <= 12'hb27;
      20'h05c7d: out <= 12'hee9;
      20'h05c7e: out <= 12'hee9;
      20'h05c7f: out <= 12'hee9;
      20'h05c80: out <= 12'h000;
      20'h05c81: out <= 12'h000;
      20'h05c82: out <= 12'h000;
      20'h05c83: out <= 12'h000;
      20'h05c84: out <= 12'h000;
      20'h05c85: out <= 12'h000;
      20'h05c86: out <= 12'h000;
      20'h05c87: out <= 12'h000;
      20'h05c88: out <= 12'h000;
      20'h05c89: out <= 12'h000;
      20'h05c8a: out <= 12'h000;
      20'h05c8b: out <= 12'h000;
      20'h05c8c: out <= 12'h603;
      20'h05c8d: out <= 12'h603;
      20'h05c8e: out <= 12'h603;
      20'h05c8f: out <= 12'h603;
      20'h05c90: out <= 12'h603;
      20'h05c91: out <= 12'h603;
      20'h05c92: out <= 12'h603;
      20'h05c93: out <= 12'h603;
      20'h05c94: out <= 12'hfff;
      20'h05c95: out <= 12'hbbb;
      20'h05c96: out <= 12'h666;
      20'h05c97: out <= 12'hfff;
      20'h05c98: out <= 12'hfff;
      20'h05c99: out <= 12'hbbb;
      20'h05c9a: out <= 12'h666;
      20'h05c9b: out <= 12'h666;
      20'h05c9c: out <= 12'hfff;
      20'h05c9d: out <= 12'h8d0;
      20'h05c9e: out <= 12'h8d0;
      20'h05c9f: out <= 12'h380;
      20'h05ca0: out <= 12'h8d0;
      20'h05ca1: out <= 12'h8d0;
      20'h05ca2: out <= 12'h000;
      20'h05ca3: out <= 12'h380;
      20'h05ca4: out <= 12'hfff;
      20'h05ca5: out <= 12'h666;
      20'h05ca6: out <= 12'h000;
      20'h05ca7: out <= 12'h000;
      20'h05ca8: out <= 12'hfff;
      20'h05ca9: out <= 12'h666;
      20'h05caa: out <= 12'h000;
      20'h05cab: out <= 12'h000;
      20'h05cac: out <= 12'hfff;
      20'h05cad: out <= 12'h6af;
      20'h05cae: out <= 12'h6af;
      20'h05caf: out <= 12'hfff;
      20'h05cb0: out <= 12'h4cd;
      20'h05cb1: out <= 12'h4cd;
      20'h05cb2: out <= 12'h4cd;
      20'h05cb3: out <= 12'h4cd;
      20'h05cb4: out <= 12'h603;
      20'h05cb5: out <= 12'h603;
      20'h05cb6: out <= 12'h603;
      20'h05cb7: out <= 12'h603;
      20'h05cb8: out <= 12'hee9;
      20'h05cb9: out <= 12'hf87;
      20'h05cba: out <= 12'hee9;
      20'h05cbb: out <= 12'hf87;
      20'h05cbc: out <= 12'hf87;
      20'h05cbd: out <= 12'hb27;
      20'h05cbe: out <= 12'hf87;
      20'h05cbf: out <= 12'hb27;
      20'h05cc0: out <= 12'h000;
      20'h05cc1: out <= 12'h000;
      20'h05cc2: out <= 12'h000;
      20'h05cc3: out <= 12'h000;
      20'h05cc4: out <= 12'h000;
      20'h05cc5: out <= 12'h000;
      20'h05cc6: out <= 12'h000;
      20'h05cc7: out <= 12'h000;
      20'h05cc8: out <= 12'h000;
      20'h05cc9: out <= 12'h6af;
      20'h05cca: out <= 12'hfff;
      20'h05ccb: out <= 12'h6af;
      20'h05ccc: out <= 12'h16d;
      20'h05ccd: out <= 12'hfff;
      20'h05cce: out <= 12'h6af;
      20'h05ccf: out <= 12'h6af;
      20'h05cd0: out <= 12'h6af;
      20'h05cd1: out <= 12'h6af;
      20'h05cd2: out <= 12'h6af;
      20'h05cd3: out <= 12'hfff;
      20'h05cd4: out <= 12'h16d;
      20'h05cd5: out <= 12'h6af;
      20'h05cd6: out <= 12'hfff;
      20'h05cd7: out <= 12'h6af;
      20'h05cd8: out <= 12'h000;
      20'h05cd9: out <= 12'h000;
      20'h05cda: out <= 12'h000;
      20'h05cdb: out <= 12'h4cd;
      20'h05cdc: out <= 12'h000;
      20'h05cdd: out <= 12'h4cd;
      20'h05cde: out <= 12'h000;
      20'h05cdf: out <= 12'h000;
      20'h05ce0: out <= 12'h4cd;
      20'h05ce1: out <= 12'h4cd;
      20'h05ce2: out <= 12'h4cd;
      20'h05ce3: out <= 12'h4cd;
      20'h05ce4: out <= 12'h4cd;
      20'h05ce5: out <= 12'h4cd;
      20'h05ce6: out <= 12'h4cd;
      20'h05ce7: out <= 12'h4cd;
      20'h05ce8: out <= 12'h5ef;
      20'h05ce9: out <= 12'h5ef;
      20'h05cea: out <= 12'h5ef;
      20'h05ceb: out <= 12'h5ef;
      20'h05cec: out <= 12'h5ef;
      20'h05ced: out <= 12'h5ef;
      20'h05cee: out <= 12'h5ef;
      20'h05cef: out <= 12'h5ef;
      20'h05cf0: out <= 12'h000;
      20'h05cf1: out <= 12'h000;
      20'h05cf2: out <= 12'h000;
      20'h05cf3: out <= 12'h000;
      20'h05cf4: out <= 12'h000;
      20'h05cf5: out <= 12'h000;
      20'h05cf6: out <= 12'h000;
      20'h05cf7: out <= 12'h000;
      20'h05cf8: out <= 12'h000;
      20'h05cf9: out <= 12'h666;
      20'h05cfa: out <= 12'hbbb;
      20'h05cfb: out <= 12'hfff;
      20'h05cfc: out <= 12'hfff;
      20'h05cfd: out <= 12'hfff;
      20'h05cfe: out <= 12'hfff;
      20'h05cff: out <= 12'hfff;
      20'h05d00: out <= 12'hfff;
      20'h05d01: out <= 12'hfff;
      20'h05d02: out <= 12'h666;
      20'h05d03: out <= 12'hbbb;
      20'h05d04: out <= 12'h666;
      20'h05d05: out <= 12'h000;
      20'h05d06: out <= 12'h000;
      20'h05d07: out <= 12'h000;
      20'h05d08: out <= 12'h222;
      20'h05d09: out <= 12'h666;
      20'h05d0a: out <= 12'hbbb;
      20'h05d0b: out <= 12'hfff;
      20'h05d0c: out <= 12'hfff;
      20'h05d0d: out <= 12'hfff;
      20'h05d0e: out <= 12'hfff;
      20'h05d0f: out <= 12'hfff;
      20'h05d10: out <= 12'hfff;
      20'h05d11: out <= 12'hfff;
      20'h05d12: out <= 12'h666;
      20'h05d13: out <= 12'hbbb;
      20'h05d14: out <= 12'h666;
      20'h05d15: out <= 12'h222;
      20'h05d16: out <= 12'h222;
      20'h05d17: out <= 12'h222;
      20'h05d18: out <= 12'h000;
      20'h05d19: out <= 12'h000;
      20'h05d1a: out <= 12'h000;
      20'h05d1b: out <= 12'h666;
      20'h05d1c: out <= 12'h666;
      20'h05d1d: out <= 12'hbbb;
      20'h05d1e: out <= 12'h666;
      20'h05d1f: out <= 12'h666;
      20'h05d20: out <= 12'hbbb;
      20'h05d21: out <= 12'h666;
      20'h05d22: out <= 12'h666;
      20'h05d23: out <= 12'hbbb;
      20'h05d24: out <= 12'h666;
      20'h05d25: out <= 12'hbbb;
      20'h05d26: out <= 12'h000;
      20'h05d27: out <= 12'h000;
      20'h05d28: out <= 12'h222;
      20'h05d29: out <= 12'h222;
      20'h05d2a: out <= 12'h222;
      20'h05d2b: out <= 12'hbbb;
      20'h05d2c: out <= 12'h666;
      20'h05d2d: out <= 12'hbbb;
      20'h05d2e: out <= 12'h666;
      20'h05d2f: out <= 12'h666;
      20'h05d30: out <= 12'hbbb;
      20'h05d31: out <= 12'h666;
      20'h05d32: out <= 12'h666;
      20'h05d33: out <= 12'hbbb;
      20'h05d34: out <= 12'h666;
      20'h05d35: out <= 12'h666;
      20'h05d36: out <= 12'h222;
      20'h05d37: out <= 12'h222;
      20'h05d38: out <= 12'h000;
      20'h05d39: out <= 12'h000;
      20'h05d3a: out <= 12'h000;
      20'h05d3b: out <= 12'h666;
      20'h05d3c: out <= 12'hbbb;
      20'h05d3d: out <= 12'h666;
      20'h05d3e: out <= 12'hfff;
      20'h05d3f: out <= 12'hfff;
      20'h05d40: out <= 12'hfff;
      20'h05d41: out <= 12'hfff;
      20'h05d42: out <= 12'hfff;
      20'h05d43: out <= 12'hfff;
      20'h05d44: out <= 12'hfff;
      20'h05d45: out <= 12'hbbb;
      20'h05d46: out <= 12'h666;
      20'h05d47: out <= 12'h000;
      20'h05d48: out <= 12'h222;
      20'h05d49: out <= 12'h222;
      20'h05d4a: out <= 12'h222;
      20'h05d4b: out <= 12'h666;
      20'h05d4c: out <= 12'hbbb;
      20'h05d4d: out <= 12'h666;
      20'h05d4e: out <= 12'hfff;
      20'h05d4f: out <= 12'hfff;
      20'h05d50: out <= 12'hfff;
      20'h05d51: out <= 12'hfff;
      20'h05d52: out <= 12'hfff;
      20'h05d53: out <= 12'hfff;
      20'h05d54: out <= 12'hfff;
      20'h05d55: out <= 12'hbbb;
      20'h05d56: out <= 12'h666;
      20'h05d57: out <= 12'h222;
      20'h05d58: out <= 12'h000;
      20'h05d59: out <= 12'h000;
      20'h05d5a: out <= 12'h000;
      20'h05d5b: out <= 12'hbbb;
      20'h05d5c: out <= 12'h666;
      20'h05d5d: out <= 12'hbbb;
      20'h05d5e: out <= 12'hfff;
      20'h05d5f: out <= 12'h666;
      20'h05d60: out <= 12'hfff;
      20'h05d61: out <= 12'hfff;
      20'h05d62: out <= 12'h666;
      20'h05d63: out <= 12'hbbb;
      20'h05d64: out <= 12'h666;
      20'h05d65: out <= 12'h666;
      20'h05d66: out <= 12'h000;
      20'h05d67: out <= 12'h000;
      20'h05d68: out <= 12'h222;
      20'h05d69: out <= 12'h222;
      20'h05d6a: out <= 12'h222;
      20'h05d6b: out <= 12'h666;
      20'h05d6c: out <= 12'h666;
      20'h05d6d: out <= 12'hbbb;
      20'h05d6e: out <= 12'hfff;
      20'h05d6f: out <= 12'h666;
      20'h05d70: out <= 12'hfff;
      20'h05d71: out <= 12'hfff;
      20'h05d72: out <= 12'h666;
      20'h05d73: out <= 12'hbbb;
      20'h05d74: out <= 12'h666;
      20'h05d75: out <= 12'hbbb;
      20'h05d76: out <= 12'h222;
      20'h05d77: out <= 12'h222;
      20'h05d78: out <= 12'h603;
      20'h05d79: out <= 12'h603;
      20'h05d7a: out <= 12'h603;
      20'h05d7b: out <= 12'h603;
      20'h05d7c: out <= 12'hb27;
      20'h05d7d: out <= 12'hf87;
      20'h05d7e: out <= 12'hf87;
      20'h05d7f: out <= 12'hf87;
      20'h05d80: out <= 12'hf87;
      20'h05d81: out <= 12'hf87;
      20'h05d82: out <= 12'hf87;
      20'h05d83: out <= 12'hee9;
      20'h05d84: out <= 12'h000;
      20'h05d85: out <= 12'h000;
      20'h05d86: out <= 12'h000;
      20'h05d87: out <= 12'h000;
      20'h05d88: out <= 12'hf87;
      20'h05d89: out <= 12'hf87;
      20'h05d8a: out <= 12'hf87;
      20'h05d8b: out <= 12'hee9;
      20'h05d8c: out <= 12'hb27;
      20'h05d8d: out <= 12'hf87;
      20'h05d8e: out <= 12'hf87;
      20'h05d8f: out <= 12'hf87;
      20'h05d90: out <= 12'hf87;
      20'h05d91: out <= 12'hf87;
      20'h05d92: out <= 12'hf87;
      20'h05d93: out <= 12'hee9;
      20'h05d94: out <= 12'hb27;
      20'h05d95: out <= 12'hf87;
      20'h05d96: out <= 12'hf87;
      20'h05d97: out <= 12'hf87;
      20'h05d98: out <= 12'h000;
      20'h05d99: out <= 12'h000;
      20'h05d9a: out <= 12'h000;
      20'h05d9b: out <= 12'h000;
      20'h05d9c: out <= 12'h000;
      20'h05d9d: out <= 12'h000;
      20'h05d9e: out <= 12'h000;
      20'h05d9f: out <= 12'h000;
      20'h05da0: out <= 12'h000;
      20'h05da1: out <= 12'h000;
      20'h05da2: out <= 12'h000;
      20'h05da3: out <= 12'h000;
      20'h05da4: out <= 12'h603;
      20'h05da5: out <= 12'h603;
      20'h05da6: out <= 12'h603;
      20'h05da7: out <= 12'h603;
      20'h05da8: out <= 12'h603;
      20'h05da9: out <= 12'h603;
      20'h05daa: out <= 12'h603;
      20'h05dab: out <= 12'h603;
      20'h05dac: out <= 12'hfff;
      20'h05dad: out <= 12'hbbb;
      20'h05dae: out <= 12'hbbb;
      20'h05daf: out <= 12'hbbb;
      20'h05db0: out <= 12'hbbb;
      20'h05db1: out <= 12'hbbb;
      20'h05db2: out <= 12'h666;
      20'h05db3: out <= 12'h666;
      20'h05db4: out <= 12'h380;
      20'h05db5: out <= 12'h8d0;
      20'h05db6: out <= 12'h380;
      20'h05db7: out <= 12'h380;
      20'h05db8: out <= 12'h8d0;
      20'h05db9: out <= 12'h380;
      20'h05dba: out <= 12'h380;
      20'h05dbb: out <= 12'h380;
      20'h05dbc: out <= 12'hbbb;
      20'h05dbd: out <= 12'hfff;
      20'h05dbe: out <= 12'h000;
      20'h05dbf: out <= 12'h000;
      20'h05dc0: out <= 12'hbbb;
      20'h05dc1: out <= 12'hfff;
      20'h05dc2: out <= 12'h000;
      20'h05dc3: out <= 12'h000;
      20'h05dc4: out <= 12'h4cd;
      20'h05dc5: out <= 12'hfff;
      20'h05dc6: out <= 12'hfff;
      20'h05dc7: out <= 12'h4cd;
      20'h05dc8: out <= 12'h4cd;
      20'h05dc9: out <= 12'h6af;
      20'h05dca: out <= 12'h6af;
      20'h05dcb: out <= 12'h4cd;
      20'h05dcc: out <= 12'h603;
      20'h05dcd: out <= 12'h603;
      20'h05dce: out <= 12'h603;
      20'h05dcf: out <= 12'h603;
      20'h05dd0: out <= 12'hee9;
      20'h05dd1: out <= 12'hf87;
      20'h05dd2: out <= 12'hee9;
      20'h05dd3: out <= 12'hb27;
      20'h05dd4: out <= 12'hb27;
      20'h05dd5: out <= 12'hb27;
      20'h05dd6: out <= 12'hf87;
      20'h05dd7: out <= 12'hb27;
      20'h05dd8: out <= 12'h000;
      20'h05dd9: out <= 12'h000;
      20'h05dda: out <= 12'h000;
      20'h05ddb: out <= 12'h000;
      20'h05ddc: out <= 12'h000;
      20'h05ddd: out <= 12'h000;
      20'h05dde: out <= 12'h000;
      20'h05ddf: out <= 12'h000;
      20'h05de0: out <= 12'h000;
      20'h05de1: out <= 12'h6af;
      20'h05de2: out <= 12'h16d;
      20'h05de3: out <= 12'h6af;
      20'h05de4: out <= 12'h000;
      20'h05de5: out <= 12'h16d;
      20'h05de6: out <= 12'h16d;
      20'h05de7: out <= 12'h16d;
      20'h05de8: out <= 12'h16d;
      20'h05de9: out <= 12'h16d;
      20'h05dea: out <= 12'h16d;
      20'h05deb: out <= 12'h16d;
      20'h05dec: out <= 12'h000;
      20'h05ded: out <= 12'h6af;
      20'h05dee: out <= 12'h16d;
      20'h05def: out <= 12'h6af;
      20'h05df0: out <= 12'h000;
      20'h05df1: out <= 12'h000;
      20'h05df2: out <= 12'h4cd;
      20'h05df3: out <= 12'h000;
      20'h05df4: out <= 12'h000;
      20'h05df5: out <= 12'h000;
      20'h05df6: out <= 12'h4cd;
      20'h05df7: out <= 12'h000;
      20'h05df8: out <= 12'h4cd;
      20'h05df9: out <= 12'h4cd;
      20'h05dfa: out <= 12'h4cd;
      20'h05dfb: out <= 12'h4cd;
      20'h05dfc: out <= 12'h4cd;
      20'h05dfd: out <= 12'h4cd;
      20'h05dfe: out <= 12'h4cd;
      20'h05dff: out <= 12'h4cd;
      20'h05e00: out <= 12'h5ef;
      20'h05e01: out <= 12'h5ef;
      20'h05e02: out <= 12'h5ef;
      20'h05e03: out <= 12'h5ef;
      20'h05e04: out <= 12'h5ef;
      20'h05e05: out <= 12'h5ef;
      20'h05e06: out <= 12'h5ef;
      20'h05e07: out <= 12'h5ef;
      20'h05e08: out <= 12'h000;
      20'h05e09: out <= 12'h000;
      20'h05e0a: out <= 12'h000;
      20'h05e0b: out <= 12'h000;
      20'h05e0c: out <= 12'h000;
      20'h05e0d: out <= 12'h000;
      20'h05e0e: out <= 12'h000;
      20'h05e0f: out <= 12'h000;
      20'h05e10: out <= 12'h000;
      20'h05e11: out <= 12'h666;
      20'h05e12: out <= 12'hbbb;
      20'h05e13: out <= 12'h666;
      20'h05e14: out <= 12'hbbb;
      20'h05e15: out <= 12'h666;
      20'h05e16: out <= 12'h666;
      20'h05e17: out <= 12'h666;
      20'h05e18: out <= 12'hbbb;
      20'h05e19: out <= 12'hfff;
      20'h05e1a: out <= 12'h666;
      20'h05e1b: out <= 12'h666;
      20'h05e1c: out <= 12'h666;
      20'h05e1d: out <= 12'h666;
      20'h05e1e: out <= 12'h666;
      20'h05e1f: out <= 12'h666;
      20'h05e20: out <= 12'h222;
      20'h05e21: out <= 12'h666;
      20'h05e22: out <= 12'hbbb;
      20'h05e23: out <= 12'h666;
      20'h05e24: out <= 12'hbbb;
      20'h05e25: out <= 12'h666;
      20'h05e26: out <= 12'h666;
      20'h05e27: out <= 12'h666;
      20'h05e28: out <= 12'hbbb;
      20'h05e29: out <= 12'hfff;
      20'h05e2a: out <= 12'h666;
      20'h05e2b: out <= 12'h666;
      20'h05e2c: out <= 12'h666;
      20'h05e2d: out <= 12'h666;
      20'h05e2e: out <= 12'h666;
      20'h05e2f: out <= 12'h666;
      20'h05e30: out <= 12'h000;
      20'h05e31: out <= 12'h000;
      20'h05e32: out <= 12'h000;
      20'h05e33: out <= 12'hbbb;
      20'h05e34: out <= 12'h666;
      20'h05e35: out <= 12'h666;
      20'h05e36: out <= 12'hfff;
      20'h05e37: out <= 12'hfff;
      20'h05e38: out <= 12'hfff;
      20'h05e39: out <= 12'hfff;
      20'h05e3a: out <= 12'hfff;
      20'h05e3b: out <= 12'h666;
      20'h05e3c: out <= 12'h666;
      20'h05e3d: out <= 12'h666;
      20'h05e3e: out <= 12'h000;
      20'h05e3f: out <= 12'h000;
      20'h05e40: out <= 12'h222;
      20'h05e41: out <= 12'h222;
      20'h05e42: out <= 12'h222;
      20'h05e43: out <= 12'h666;
      20'h05e44: out <= 12'h666;
      20'h05e45: out <= 12'h666;
      20'h05e46: out <= 12'hfff;
      20'h05e47: out <= 12'hfff;
      20'h05e48: out <= 12'hfff;
      20'h05e49: out <= 12'hfff;
      20'h05e4a: out <= 12'hfff;
      20'h05e4b: out <= 12'h666;
      20'h05e4c: out <= 12'h666;
      20'h05e4d: out <= 12'hbbb;
      20'h05e4e: out <= 12'h222;
      20'h05e4f: out <= 12'h222;
      20'h05e50: out <= 12'h666;
      20'h05e51: out <= 12'h666;
      20'h05e52: out <= 12'h666;
      20'h05e53: out <= 12'h666;
      20'h05e54: out <= 12'h666;
      20'h05e55: out <= 12'h666;
      20'h05e56: out <= 12'hfff;
      20'h05e57: out <= 12'hbbb;
      20'h05e58: out <= 12'h666;
      20'h05e59: out <= 12'h666;
      20'h05e5a: out <= 12'h666;
      20'h05e5b: out <= 12'hbbb;
      20'h05e5c: out <= 12'h666;
      20'h05e5d: out <= 12'hbbb;
      20'h05e5e: out <= 12'h666;
      20'h05e5f: out <= 12'h000;
      20'h05e60: out <= 12'h666;
      20'h05e61: out <= 12'h666;
      20'h05e62: out <= 12'h666;
      20'h05e63: out <= 12'h666;
      20'h05e64: out <= 12'h666;
      20'h05e65: out <= 12'h666;
      20'h05e66: out <= 12'hfff;
      20'h05e67: out <= 12'hbbb;
      20'h05e68: out <= 12'h666;
      20'h05e69: out <= 12'h666;
      20'h05e6a: out <= 12'h666;
      20'h05e6b: out <= 12'hbbb;
      20'h05e6c: out <= 12'h666;
      20'h05e6d: out <= 12'hbbb;
      20'h05e6e: out <= 12'h666;
      20'h05e6f: out <= 12'h222;
      20'h05e70: out <= 12'h000;
      20'h05e71: out <= 12'h000;
      20'h05e72: out <= 12'h000;
      20'h05e73: out <= 12'h666;
      20'h05e74: out <= 12'h666;
      20'h05e75: out <= 12'hbbb;
      20'h05e76: out <= 12'hfff;
      20'h05e77: out <= 12'h666;
      20'h05e78: out <= 12'hbbb;
      20'h05e79: out <= 12'hfff;
      20'h05e7a: out <= 12'h666;
      20'h05e7b: out <= 12'hbbb;
      20'h05e7c: out <= 12'h666;
      20'h05e7d: out <= 12'hbbb;
      20'h05e7e: out <= 12'h000;
      20'h05e7f: out <= 12'h000;
      20'h05e80: out <= 12'h222;
      20'h05e81: out <= 12'h222;
      20'h05e82: out <= 12'h222;
      20'h05e83: out <= 12'hbbb;
      20'h05e84: out <= 12'h666;
      20'h05e85: out <= 12'hbbb;
      20'h05e86: out <= 12'hfff;
      20'h05e87: out <= 12'h666;
      20'h05e88: out <= 12'hbbb;
      20'h05e89: out <= 12'hfff;
      20'h05e8a: out <= 12'h666;
      20'h05e8b: out <= 12'hbbb;
      20'h05e8c: out <= 12'h666;
      20'h05e8d: out <= 12'h666;
      20'h05e8e: out <= 12'h222;
      20'h05e8f: out <= 12'h222;
      20'h05e90: out <= 12'h603;
      20'h05e91: out <= 12'h603;
      20'h05e92: out <= 12'h603;
      20'h05e93: out <= 12'h603;
      20'h05e94: out <= 12'hb27;
      20'h05e95: out <= 12'hf87;
      20'h05e96: out <= 12'hf87;
      20'h05e97: out <= 12'hf87;
      20'h05e98: out <= 12'hf87;
      20'h05e99: out <= 12'hf87;
      20'h05e9a: out <= 12'hf87;
      20'h05e9b: out <= 12'hee9;
      20'h05e9c: out <= 12'h000;
      20'h05e9d: out <= 12'h000;
      20'h05e9e: out <= 12'h000;
      20'h05e9f: out <= 12'h000;
      20'h05ea0: out <= 12'hf87;
      20'h05ea1: out <= 12'hf87;
      20'h05ea2: out <= 12'hf87;
      20'h05ea3: out <= 12'hee9;
      20'h05ea4: out <= 12'hb27;
      20'h05ea5: out <= 12'hf87;
      20'h05ea6: out <= 12'hf87;
      20'h05ea7: out <= 12'hf87;
      20'h05ea8: out <= 12'hf87;
      20'h05ea9: out <= 12'hf87;
      20'h05eaa: out <= 12'hf87;
      20'h05eab: out <= 12'hee9;
      20'h05eac: out <= 12'hb27;
      20'h05ead: out <= 12'hf87;
      20'h05eae: out <= 12'hf87;
      20'h05eaf: out <= 12'hf87;
      20'h05eb0: out <= 12'h000;
      20'h05eb1: out <= 12'h000;
      20'h05eb2: out <= 12'h000;
      20'h05eb3: out <= 12'h000;
      20'h05eb4: out <= 12'h000;
      20'h05eb5: out <= 12'h000;
      20'h05eb6: out <= 12'h000;
      20'h05eb7: out <= 12'h000;
      20'h05eb8: out <= 12'h000;
      20'h05eb9: out <= 12'h000;
      20'h05eba: out <= 12'h000;
      20'h05ebb: out <= 12'h000;
      20'h05ebc: out <= 12'h603;
      20'h05ebd: out <= 12'h603;
      20'h05ebe: out <= 12'h603;
      20'h05ebf: out <= 12'h603;
      20'h05ec0: out <= 12'h603;
      20'h05ec1: out <= 12'h603;
      20'h05ec2: out <= 12'h603;
      20'h05ec3: out <= 12'h603;
      20'h05ec4: out <= 12'hfff;
      20'h05ec5: out <= 12'h666;
      20'h05ec6: out <= 12'h666;
      20'h05ec7: out <= 12'h666;
      20'h05ec8: out <= 12'h666;
      20'h05ec9: out <= 12'h666;
      20'h05eca: out <= 12'h666;
      20'h05ecb: out <= 12'h666;
      20'h05ecc: out <= 12'h000;
      20'h05ecd: out <= 12'h380;
      20'h05ece: out <= 12'h8d0;
      20'h05ecf: out <= 12'h8d0;
      20'h05ed0: out <= 12'h000;
      20'h05ed1: out <= 12'h380;
      20'h05ed2: out <= 12'h000;
      20'h05ed3: out <= 12'h380;
      20'h05ed4: out <= 12'h000;
      20'h05ed5: out <= 12'h000;
      20'h05ed6: out <= 12'hfff;
      20'h05ed7: out <= 12'h666;
      20'h05ed8: out <= 12'h000;
      20'h05ed9: out <= 12'h000;
      20'h05eda: out <= 12'hfff;
      20'h05edb: out <= 12'h666;
      20'h05edc: out <= 12'h4cd;
      20'h05edd: out <= 12'h4cd;
      20'h05ede: out <= 12'h4cd;
      20'h05edf: out <= 12'h4cd;
      20'h05ee0: out <= 12'h6af;
      20'h05ee1: out <= 12'hfff;
      20'h05ee2: out <= 12'hfff;
      20'h05ee3: out <= 12'h6af;
      20'h05ee4: out <= 12'h603;
      20'h05ee5: out <= 12'h603;
      20'h05ee6: out <= 12'h603;
      20'h05ee7: out <= 12'h603;
      20'h05ee8: out <= 12'hee9;
      20'h05ee9: out <= 12'hf87;
      20'h05eea: out <= 12'hf87;
      20'h05eeb: out <= 12'hf87;
      20'h05eec: out <= 12'hf87;
      20'h05eed: out <= 12'hf87;
      20'h05eee: out <= 12'hf87;
      20'h05eef: out <= 12'hb27;
      20'h05ef0: out <= 12'h000;
      20'h05ef1: out <= 12'h000;
      20'h05ef2: out <= 12'h000;
      20'h05ef3: out <= 12'h000;
      20'h05ef4: out <= 12'h000;
      20'h05ef5: out <= 12'h000;
      20'h05ef6: out <= 12'h000;
      20'h05ef7: out <= 12'h000;
      20'h05ef8: out <= 12'h000;
      20'h05ef9: out <= 12'h6af;
      20'h05efa: out <= 12'hfff;
      20'h05efb: out <= 12'h6af;
      20'h05efc: out <= 12'h000;
      20'h05efd: out <= 12'h000;
      20'h05efe: out <= 12'h000;
      20'h05eff: out <= 12'h000;
      20'h05f00: out <= 12'h000;
      20'h05f01: out <= 12'h000;
      20'h05f02: out <= 12'h000;
      20'h05f03: out <= 12'h000;
      20'h05f04: out <= 12'h000;
      20'h05f05: out <= 12'h6af;
      20'h05f06: out <= 12'hfff;
      20'h05f07: out <= 12'h6af;
      20'h05f08: out <= 12'h000;
      20'h05f09: out <= 12'h000;
      20'h05f0a: out <= 12'h000;
      20'h05f0b: out <= 12'h000;
      20'h05f0c: out <= 12'h000;
      20'h05f0d: out <= 12'h000;
      20'h05f0e: out <= 12'h000;
      20'h05f0f: out <= 12'h000;
      20'h05f10: out <= 12'h4cd;
      20'h05f11: out <= 12'h4cd;
      20'h05f12: out <= 12'h4cd;
      20'h05f13: out <= 12'h4cd;
      20'h05f14: out <= 12'h4cd;
      20'h05f15: out <= 12'h4cd;
      20'h05f16: out <= 12'h4cd;
      20'h05f17: out <= 12'h4cd;
      20'h05f18: out <= 12'h5ef;
      20'h05f19: out <= 12'h5ef;
      20'h05f1a: out <= 12'h5ef;
      20'h05f1b: out <= 12'h5ef;
      20'h05f1c: out <= 12'h5ef;
      20'h05f1d: out <= 12'h5ef;
      20'h05f1e: out <= 12'h5ef;
      20'h05f1f: out <= 12'h5ef;
      20'h05f20: out <= 12'h000;
      20'h05f21: out <= 12'h000;
      20'h05f22: out <= 12'h000;
      20'h05f23: out <= 12'h000;
      20'h05f24: out <= 12'h000;
      20'h05f25: out <= 12'h000;
      20'h05f26: out <= 12'h000;
      20'h05f27: out <= 12'h000;
      20'h05f28: out <= 12'h000;
      20'h05f29: out <= 12'h666;
      20'h05f2a: out <= 12'hbbb;
      20'h05f2b: out <= 12'h666;
      20'h05f2c: out <= 12'hbbb;
      20'h05f2d: out <= 12'hfff;
      20'h05f2e: out <= 12'hbbb;
      20'h05f2f: out <= 12'h666;
      20'h05f30: out <= 12'hbbb;
      20'h05f31: out <= 12'hfff;
      20'h05f32: out <= 12'hbbb;
      20'h05f33: out <= 12'hbbb;
      20'h05f34: out <= 12'hfff;
      20'h05f35: out <= 12'hfff;
      20'h05f36: out <= 12'hfff;
      20'h05f37: out <= 12'hfff;
      20'h05f38: out <= 12'h222;
      20'h05f39: out <= 12'h666;
      20'h05f3a: out <= 12'hbbb;
      20'h05f3b: out <= 12'h666;
      20'h05f3c: out <= 12'hbbb;
      20'h05f3d: out <= 12'hfff;
      20'h05f3e: out <= 12'hbbb;
      20'h05f3f: out <= 12'h666;
      20'h05f40: out <= 12'hbbb;
      20'h05f41: out <= 12'hfff;
      20'h05f42: out <= 12'hbbb;
      20'h05f43: out <= 12'hbbb;
      20'h05f44: out <= 12'hfff;
      20'h05f45: out <= 12'hfff;
      20'h05f46: out <= 12'hfff;
      20'h05f47: out <= 12'hfff;
      20'h05f48: out <= 12'h000;
      20'h05f49: out <= 12'h000;
      20'h05f4a: out <= 12'h000;
      20'h05f4b: out <= 12'h666;
      20'h05f4c: out <= 12'h666;
      20'h05f4d: out <= 12'hbbb;
      20'h05f4e: out <= 12'hfff;
      20'h05f4f: out <= 12'hbbb;
      20'h05f50: out <= 12'hbbb;
      20'h05f51: out <= 12'hbbb;
      20'h05f52: out <= 12'h666;
      20'h05f53: out <= 12'hbbb;
      20'h05f54: out <= 12'h666;
      20'h05f55: out <= 12'hbbb;
      20'h05f56: out <= 12'h000;
      20'h05f57: out <= 12'h000;
      20'h05f58: out <= 12'h222;
      20'h05f59: out <= 12'h222;
      20'h05f5a: out <= 12'h222;
      20'h05f5b: out <= 12'hbbb;
      20'h05f5c: out <= 12'h666;
      20'h05f5d: out <= 12'hbbb;
      20'h05f5e: out <= 12'hfff;
      20'h05f5f: out <= 12'hbbb;
      20'h05f60: out <= 12'hbbb;
      20'h05f61: out <= 12'hbbb;
      20'h05f62: out <= 12'h666;
      20'h05f63: out <= 12'hbbb;
      20'h05f64: out <= 12'h666;
      20'h05f65: out <= 12'h666;
      20'h05f66: out <= 12'h222;
      20'h05f67: out <= 12'h222;
      20'h05f68: out <= 12'hfff;
      20'h05f69: out <= 12'hfff;
      20'h05f6a: out <= 12'hfff;
      20'h05f6b: out <= 12'hfff;
      20'h05f6c: out <= 12'hbbb;
      20'h05f6d: out <= 12'hbbb;
      20'h05f6e: out <= 12'hfff;
      20'h05f6f: out <= 12'hbbb;
      20'h05f70: out <= 12'h666;
      20'h05f71: out <= 12'hbbb;
      20'h05f72: out <= 12'hfff;
      20'h05f73: out <= 12'hbbb;
      20'h05f74: out <= 12'h666;
      20'h05f75: out <= 12'hbbb;
      20'h05f76: out <= 12'h666;
      20'h05f77: out <= 12'h000;
      20'h05f78: out <= 12'hfff;
      20'h05f79: out <= 12'hfff;
      20'h05f7a: out <= 12'hfff;
      20'h05f7b: out <= 12'hfff;
      20'h05f7c: out <= 12'hbbb;
      20'h05f7d: out <= 12'hbbb;
      20'h05f7e: out <= 12'hfff;
      20'h05f7f: out <= 12'hbbb;
      20'h05f80: out <= 12'h666;
      20'h05f81: out <= 12'hbbb;
      20'h05f82: out <= 12'hfff;
      20'h05f83: out <= 12'hbbb;
      20'h05f84: out <= 12'h666;
      20'h05f85: out <= 12'hbbb;
      20'h05f86: out <= 12'h666;
      20'h05f87: out <= 12'h222;
      20'h05f88: out <= 12'h000;
      20'h05f89: out <= 12'h000;
      20'h05f8a: out <= 12'h000;
      20'h05f8b: out <= 12'hbbb;
      20'h05f8c: out <= 12'h666;
      20'h05f8d: out <= 12'hbbb;
      20'h05f8e: out <= 12'hfff;
      20'h05f8f: out <= 12'h666;
      20'h05f90: out <= 12'h666;
      20'h05f91: out <= 12'h666;
      20'h05f92: out <= 12'h666;
      20'h05f93: out <= 12'hbbb;
      20'h05f94: out <= 12'h666;
      20'h05f95: out <= 12'h666;
      20'h05f96: out <= 12'h000;
      20'h05f97: out <= 12'h000;
      20'h05f98: out <= 12'h222;
      20'h05f99: out <= 12'h222;
      20'h05f9a: out <= 12'h222;
      20'h05f9b: out <= 12'h666;
      20'h05f9c: out <= 12'h666;
      20'h05f9d: out <= 12'hbbb;
      20'h05f9e: out <= 12'hfff;
      20'h05f9f: out <= 12'h666;
      20'h05fa0: out <= 12'h666;
      20'h05fa1: out <= 12'h666;
      20'h05fa2: out <= 12'h666;
      20'h05fa3: out <= 12'hbbb;
      20'h05fa4: out <= 12'h666;
      20'h05fa5: out <= 12'hbbb;
      20'h05fa6: out <= 12'h222;
      20'h05fa7: out <= 12'h222;
      20'h05fa8: out <= 12'h603;
      20'h05fa9: out <= 12'h603;
      20'h05faa: out <= 12'h603;
      20'h05fab: out <= 12'h603;
      20'h05fac: out <= 12'hb27;
      20'h05fad: out <= 12'hb27;
      20'h05fae: out <= 12'hb27;
      20'h05faf: out <= 12'hb27;
      20'h05fb0: out <= 12'hb27;
      20'h05fb1: out <= 12'hb27;
      20'h05fb2: out <= 12'hb27;
      20'h05fb3: out <= 12'hb27;
      20'h05fb4: out <= 12'h000;
      20'h05fb5: out <= 12'h000;
      20'h05fb6: out <= 12'h000;
      20'h05fb7: out <= 12'h000;
      20'h05fb8: out <= 12'hb27;
      20'h05fb9: out <= 12'hb27;
      20'h05fba: out <= 12'hb27;
      20'h05fbb: out <= 12'hb27;
      20'h05fbc: out <= 12'hb27;
      20'h05fbd: out <= 12'hb27;
      20'h05fbe: out <= 12'hb27;
      20'h05fbf: out <= 12'hb27;
      20'h05fc0: out <= 12'hb27;
      20'h05fc1: out <= 12'hb27;
      20'h05fc2: out <= 12'hb27;
      20'h05fc3: out <= 12'hb27;
      20'h05fc4: out <= 12'hb27;
      20'h05fc5: out <= 12'hb27;
      20'h05fc6: out <= 12'hb27;
      20'h05fc7: out <= 12'hb27;
      20'h05fc8: out <= 12'h000;
      20'h05fc9: out <= 12'h000;
      20'h05fca: out <= 12'h000;
      20'h05fcb: out <= 12'h000;
      20'h05fcc: out <= 12'h000;
      20'h05fcd: out <= 12'h000;
      20'h05fce: out <= 12'h000;
      20'h05fcf: out <= 12'h000;
      20'h05fd0: out <= 12'h000;
      20'h05fd1: out <= 12'h000;
      20'h05fd2: out <= 12'h000;
      20'h05fd3: out <= 12'h000;
      20'h05fd4: out <= 12'h603;
      20'h05fd5: out <= 12'h603;
      20'h05fd6: out <= 12'h603;
      20'h05fd7: out <= 12'h603;
      20'h05fd8: out <= 12'h603;
      20'h05fd9: out <= 12'h603;
      20'h05fda: out <= 12'h603;
      20'h05fdb: out <= 12'h603;
      20'h05fdc: out <= 12'h666;
      20'h05fdd: out <= 12'h666;
      20'h05fde: out <= 12'h666;
      20'h05fdf: out <= 12'h666;
      20'h05fe0: out <= 12'h666;
      20'h05fe1: out <= 12'h666;
      20'h05fe2: out <= 12'h666;
      20'h05fe3: out <= 12'h666;
      20'h05fe4: out <= 12'h000;
      20'h05fe5: out <= 12'h000;
      20'h05fe6: out <= 12'h380;
      20'h05fe7: out <= 12'h380;
      20'h05fe8: out <= 12'h380;
      20'h05fe9: out <= 12'h380;
      20'h05fea: out <= 12'h000;
      20'h05feb: out <= 12'h000;
      20'h05fec: out <= 12'h000;
      20'h05fed: out <= 12'h000;
      20'h05fee: out <= 12'hbbb;
      20'h05fef: out <= 12'hfff;
      20'h05ff0: out <= 12'h000;
      20'h05ff1: out <= 12'h000;
      20'h05ff2: out <= 12'hbbb;
      20'h05ff3: out <= 12'hfff;
      20'h05ff4: out <= 12'h6af;
      20'h05ff5: out <= 12'h4cd;
      20'h05ff6: out <= 12'h4cd;
      20'h05ff7: out <= 12'h6af;
      20'h05ff8: out <= 12'hfff;
      20'h05ff9: out <= 12'h4cd;
      20'h05ffa: out <= 12'h4cd;
      20'h05ffb: out <= 12'hfff;
      20'h05ffc: out <= 12'h603;
      20'h05ffd: out <= 12'h603;
      20'h05ffe: out <= 12'h603;
      20'h05fff: out <= 12'h603;
      20'h06000: out <= 12'hb27;
      20'h06001: out <= 12'hb27;
      20'h06002: out <= 12'hb27;
      20'h06003: out <= 12'hb27;
      20'h06004: out <= 12'hb27;
      20'h06005: out <= 12'hb27;
      20'h06006: out <= 12'hb27;
      20'h06007: out <= 12'hb27;
      20'h06008: out <= 12'h000;
      20'h06009: out <= 12'h000;
      20'h0600a: out <= 12'h000;
      20'h0600b: out <= 12'h000;
      20'h0600c: out <= 12'h000;
      20'h0600d: out <= 12'h000;
      20'h0600e: out <= 12'h000;
      20'h0600f: out <= 12'h000;
      20'h06010: out <= 12'h000;
      20'h06011: out <= 12'h000;
      20'h06012: out <= 12'h000;
      20'h06013: out <= 12'h000;
      20'h06014: out <= 12'h000;
      20'h06015: out <= 12'h000;
      20'h06016: out <= 12'h000;
      20'h06017: out <= 12'h000;
      20'h06018: out <= 12'h000;
      20'h06019: out <= 12'h000;
      20'h0601a: out <= 12'h000;
      20'h0601b: out <= 12'h000;
      20'h0601c: out <= 12'h000;
      20'h0601d: out <= 12'h000;
      20'h0601e: out <= 12'h000;
      20'h0601f: out <= 12'h000;
      20'h06020: out <= 12'h000;
      20'h06021: out <= 12'h000;
      20'h06022: out <= 12'h000;
      20'h06023: out <= 12'h000;
      20'h06024: out <= 12'h000;
      20'h06025: out <= 12'h000;
      20'h06026: out <= 12'h000;
      20'h06027: out <= 12'h000;
      20'h06028: out <= 12'h4cd;
      20'h06029: out <= 12'h4cd;
      20'h0602a: out <= 12'h4cd;
      20'h0602b: out <= 12'h4cd;
      20'h0602c: out <= 12'h4cd;
      20'h0602d: out <= 12'h4cd;
      20'h0602e: out <= 12'h4cd;
      20'h0602f: out <= 12'h4cd;
      20'h06030: out <= 12'h5ef;
      20'h06031: out <= 12'h5ef;
      20'h06032: out <= 12'h5ef;
      20'h06033: out <= 12'h5ef;
      20'h06034: out <= 12'h5ef;
      20'h06035: out <= 12'h5ef;
      20'h06036: out <= 12'h5ef;
      20'h06037: out <= 12'h5ef;
      20'h06038: out <= 12'h000;
      20'h06039: out <= 12'h000;
      20'h0603a: out <= 12'h000;
      20'h0603b: out <= 12'h000;
      20'h0603c: out <= 12'h000;
      20'h0603d: out <= 12'h000;
      20'h0603e: out <= 12'h000;
      20'h0603f: out <= 12'h000;
      20'h06040: out <= 12'h000;
      20'h06041: out <= 12'h666;
      20'h06042: out <= 12'hbbb;
      20'h06043: out <= 12'h666;
      20'h06044: out <= 12'hbbb;
      20'h06045: out <= 12'hfff;
      20'h06046: out <= 12'hfff;
      20'h06047: out <= 12'h666;
      20'h06048: out <= 12'hbbb;
      20'h06049: out <= 12'hfff;
      20'h0604a: out <= 12'h666;
      20'h0604b: out <= 12'h666;
      20'h0604c: out <= 12'h666;
      20'h0604d: out <= 12'h666;
      20'h0604e: out <= 12'h666;
      20'h0604f: out <= 12'h666;
      20'h06050: out <= 12'h222;
      20'h06051: out <= 12'h666;
      20'h06052: out <= 12'hbbb;
      20'h06053: out <= 12'h666;
      20'h06054: out <= 12'hbbb;
      20'h06055: out <= 12'hfff;
      20'h06056: out <= 12'hfff;
      20'h06057: out <= 12'h666;
      20'h06058: out <= 12'hbbb;
      20'h06059: out <= 12'hfff;
      20'h0605a: out <= 12'h666;
      20'h0605b: out <= 12'h666;
      20'h0605c: out <= 12'h666;
      20'h0605d: out <= 12'h666;
      20'h0605e: out <= 12'h666;
      20'h0605f: out <= 12'h666;
      20'h06060: out <= 12'h000;
      20'h06061: out <= 12'h000;
      20'h06062: out <= 12'h000;
      20'h06063: out <= 12'hbbb;
      20'h06064: out <= 12'h666;
      20'h06065: out <= 12'hbbb;
      20'h06066: out <= 12'hfff;
      20'h06067: out <= 12'h666;
      20'h06068: out <= 12'h666;
      20'h06069: out <= 12'h666;
      20'h0606a: out <= 12'h666;
      20'h0606b: out <= 12'hbbb;
      20'h0606c: out <= 12'h666;
      20'h0606d: out <= 12'h666;
      20'h0606e: out <= 12'h000;
      20'h0606f: out <= 12'h000;
      20'h06070: out <= 12'h222;
      20'h06071: out <= 12'h222;
      20'h06072: out <= 12'h222;
      20'h06073: out <= 12'h666;
      20'h06074: out <= 12'h666;
      20'h06075: out <= 12'hbbb;
      20'h06076: out <= 12'hfff;
      20'h06077: out <= 12'h666;
      20'h06078: out <= 12'h666;
      20'h06079: out <= 12'h666;
      20'h0607a: out <= 12'h666;
      20'h0607b: out <= 12'hbbb;
      20'h0607c: out <= 12'h666;
      20'h0607d: out <= 12'hbbb;
      20'h0607e: out <= 12'h222;
      20'h0607f: out <= 12'h222;
      20'h06080: out <= 12'h666;
      20'h06081: out <= 12'h666;
      20'h06082: out <= 12'h666;
      20'h06083: out <= 12'h666;
      20'h06084: out <= 12'h666;
      20'h06085: out <= 12'h666;
      20'h06086: out <= 12'hfff;
      20'h06087: out <= 12'hbbb;
      20'h06088: out <= 12'h666;
      20'h06089: out <= 12'hfff;
      20'h0608a: out <= 12'hfff;
      20'h0608b: out <= 12'hbbb;
      20'h0608c: out <= 12'h666;
      20'h0608d: out <= 12'hbbb;
      20'h0608e: out <= 12'h666;
      20'h0608f: out <= 12'h000;
      20'h06090: out <= 12'h666;
      20'h06091: out <= 12'h666;
      20'h06092: out <= 12'h666;
      20'h06093: out <= 12'h666;
      20'h06094: out <= 12'h666;
      20'h06095: out <= 12'h666;
      20'h06096: out <= 12'hfff;
      20'h06097: out <= 12'hbbb;
      20'h06098: out <= 12'h666;
      20'h06099: out <= 12'hfff;
      20'h0609a: out <= 12'hfff;
      20'h0609b: out <= 12'hbbb;
      20'h0609c: out <= 12'h666;
      20'h0609d: out <= 12'hbbb;
      20'h0609e: out <= 12'h666;
      20'h0609f: out <= 12'h222;
      20'h060a0: out <= 12'h000;
      20'h060a1: out <= 12'h000;
      20'h060a2: out <= 12'h000;
      20'h060a3: out <= 12'h666;
      20'h060a4: out <= 12'h666;
      20'h060a5: out <= 12'hbbb;
      20'h060a6: out <= 12'hfff;
      20'h060a7: out <= 12'hbbb;
      20'h060a8: out <= 12'hbbb;
      20'h060a9: out <= 12'hbbb;
      20'h060aa: out <= 12'h666;
      20'h060ab: out <= 12'hbbb;
      20'h060ac: out <= 12'h666;
      20'h060ad: out <= 12'hbbb;
      20'h060ae: out <= 12'h000;
      20'h060af: out <= 12'h000;
      20'h060b0: out <= 12'h222;
      20'h060b1: out <= 12'h222;
      20'h060b2: out <= 12'h222;
      20'h060b3: out <= 12'hbbb;
      20'h060b4: out <= 12'h666;
      20'h060b5: out <= 12'hbbb;
      20'h060b6: out <= 12'hfff;
      20'h060b7: out <= 12'hbbb;
      20'h060b8: out <= 12'hbbb;
      20'h060b9: out <= 12'hbbb;
      20'h060ba: out <= 12'h666;
      20'h060bb: out <= 12'hbbb;
      20'h060bc: out <= 12'h666;
      20'h060bd: out <= 12'h666;
      20'h060be: out <= 12'h222;
      20'h060bf: out <= 12'h222;
      20'h060c0: out <= 12'h603;
      20'h060c1: out <= 12'h603;
      20'h060c2: out <= 12'h603;
      20'h060c3: out <= 12'h603;
      20'h060c4: out <= 12'h603;
      20'h060c5: out <= 12'h603;
      20'h060c6: out <= 12'h603;
      20'h060c7: out <= 12'h603;
      20'h060c8: out <= 12'h603;
      20'h060c9: out <= 12'h603;
      20'h060ca: out <= 12'h603;
      20'h060cb: out <= 12'h603;
      20'h060cc: out <= 12'h603;
      20'h060cd: out <= 12'h603;
      20'h060ce: out <= 12'h603;
      20'h060cf: out <= 12'h603;
      20'h060d0: out <= 12'h603;
      20'h060d1: out <= 12'h603;
      20'h060d2: out <= 12'h603;
      20'h060d3: out <= 12'h603;
      20'h060d4: out <= 12'h603;
      20'h060d5: out <= 12'h603;
      20'h060d6: out <= 12'h603;
      20'h060d7: out <= 12'h603;
      20'h060d8: out <= 12'h603;
      20'h060d9: out <= 12'h603;
      20'h060da: out <= 12'h603;
      20'h060db: out <= 12'h603;
      20'h060dc: out <= 12'h603;
      20'h060dd: out <= 12'h603;
      20'h060de: out <= 12'h603;
      20'h060df: out <= 12'h603;
      20'h060e0: out <= 12'h603;
      20'h060e1: out <= 12'h603;
      20'h060e2: out <= 12'h603;
      20'h060e3: out <= 12'h603;
      20'h060e4: out <= 12'h603;
      20'h060e5: out <= 12'h603;
      20'h060e6: out <= 12'h603;
      20'h060e7: out <= 12'h603;
      20'h060e8: out <= 12'h603;
      20'h060e9: out <= 12'h603;
      20'h060ea: out <= 12'h603;
      20'h060eb: out <= 12'h603;
      20'h060ec: out <= 12'h603;
      20'h060ed: out <= 12'h603;
      20'h060ee: out <= 12'h603;
      20'h060ef: out <= 12'h603;
      20'h060f0: out <= 12'h603;
      20'h060f1: out <= 12'h603;
      20'h060f2: out <= 12'h603;
      20'h060f3: out <= 12'h603;
      20'h060f4: out <= 12'h603;
      20'h060f5: out <= 12'h603;
      20'h060f6: out <= 12'h603;
      20'h060f7: out <= 12'h603;
      20'h060f8: out <= 12'h603;
      20'h060f9: out <= 12'h603;
      20'h060fa: out <= 12'h603;
      20'h060fb: out <= 12'h603;
      20'h060fc: out <= 12'h603;
      20'h060fd: out <= 12'h603;
      20'h060fe: out <= 12'h603;
      20'h060ff: out <= 12'h603;
      20'h06100: out <= 12'h603;
      20'h06101: out <= 12'h603;
      20'h06102: out <= 12'h603;
      20'h06103: out <= 12'h603;
      20'h06104: out <= 12'h603;
      20'h06105: out <= 12'h603;
      20'h06106: out <= 12'h603;
      20'h06107: out <= 12'h603;
      20'h06108: out <= 12'h603;
      20'h06109: out <= 12'h603;
      20'h0610a: out <= 12'h603;
      20'h0610b: out <= 12'h603;
      20'h0610c: out <= 12'h603;
      20'h0610d: out <= 12'h603;
      20'h0610e: out <= 12'h603;
      20'h0610f: out <= 12'h603;
      20'h06110: out <= 12'h603;
      20'h06111: out <= 12'h603;
      20'h06112: out <= 12'h603;
      20'h06113: out <= 12'h603;
      20'h06114: out <= 12'h603;
      20'h06115: out <= 12'h603;
      20'h06116: out <= 12'h603;
      20'h06117: out <= 12'h603;
      20'h06118: out <= 12'hee9;
      20'h06119: out <= 12'hee9;
      20'h0611a: out <= 12'hee9;
      20'h0611b: out <= 12'hee9;
      20'h0611c: out <= 12'hee9;
      20'h0611d: out <= 12'hee9;
      20'h0611e: out <= 12'hee9;
      20'h0611f: out <= 12'hb27;
      20'h06120: out <= 12'h000;
      20'h06121: out <= 12'h000;
      20'h06122: out <= 12'h000;
      20'h06123: out <= 12'h000;
      20'h06124: out <= 12'h000;
      20'h06125: out <= 12'h000;
      20'h06126: out <= 12'h000;
      20'h06127: out <= 12'h000;
      20'h06128: out <= 12'hfa9;
      20'h06129: out <= 12'hfa9;
      20'h0612a: out <= 12'hfa9;
      20'h0612b: out <= 12'hfa9;
      20'h0612c: out <= 12'hfa9;
      20'h0612d: out <= 12'hfa9;
      20'h0612e: out <= 12'hfa9;
      20'h0612f: out <= 12'hfa9;
      20'h06130: out <= 12'hf76;
      20'h06131: out <= 12'hf76;
      20'h06132: out <= 12'hf76;
      20'h06133: out <= 12'hf76;
      20'h06134: out <= 12'hf76;
      20'h06135: out <= 12'hf76;
      20'h06136: out <= 12'hf76;
      20'h06137: out <= 12'hf76;
      20'h06138: out <= 12'hfa9;
      20'h06139: out <= 12'hfa9;
      20'h0613a: out <= 12'hfa9;
      20'h0613b: out <= 12'hfa9;
      20'h0613c: out <= 12'hfa9;
      20'h0613d: out <= 12'hfa9;
      20'h0613e: out <= 12'hfa9;
      20'h0613f: out <= 12'hfa9;
      20'h06140: out <= 12'hf76;
      20'h06141: out <= 12'hf76;
      20'h06142: out <= 12'hf76;
      20'h06143: out <= 12'hf76;
      20'h06144: out <= 12'hf76;
      20'h06145: out <= 12'hf76;
      20'h06146: out <= 12'hf76;
      20'h06147: out <= 12'hf76;
      20'h06148: out <= 12'hfa9;
      20'h06149: out <= 12'hfa9;
      20'h0614a: out <= 12'hfa9;
      20'h0614b: out <= 12'hfa9;
      20'h0614c: out <= 12'hfa9;
      20'h0614d: out <= 12'hfa9;
      20'h0614e: out <= 12'hfa9;
      20'h0614f: out <= 12'hfa9;
      20'h06150: out <= 12'h000;
      20'h06151: out <= 12'h000;
      20'h06152: out <= 12'h000;
      20'h06153: out <= 12'h000;
      20'h06154: out <= 12'h000;
      20'h06155: out <= 12'h000;
      20'h06156: out <= 12'h000;
      20'h06157: out <= 12'h000;
      20'h06158: out <= 12'h000;
      20'h06159: out <= 12'h666;
      20'h0615a: out <= 12'hbbb;
      20'h0615b: out <= 12'h666;
      20'h0615c: out <= 12'h666;
      20'h0615d: out <= 12'h666;
      20'h0615e: out <= 12'h666;
      20'h0615f: out <= 12'h666;
      20'h06160: out <= 12'h666;
      20'h06161: out <= 12'hfff;
      20'h06162: out <= 12'h666;
      20'h06163: out <= 12'hbbb;
      20'h06164: out <= 12'h666;
      20'h06165: out <= 12'h000;
      20'h06166: out <= 12'h000;
      20'h06167: out <= 12'h000;
      20'h06168: out <= 12'h222;
      20'h06169: out <= 12'h666;
      20'h0616a: out <= 12'hbbb;
      20'h0616b: out <= 12'h666;
      20'h0616c: out <= 12'h666;
      20'h0616d: out <= 12'h666;
      20'h0616e: out <= 12'h666;
      20'h0616f: out <= 12'h666;
      20'h06170: out <= 12'h666;
      20'h06171: out <= 12'hfff;
      20'h06172: out <= 12'h666;
      20'h06173: out <= 12'hbbb;
      20'h06174: out <= 12'h666;
      20'h06175: out <= 12'h222;
      20'h06176: out <= 12'h222;
      20'h06177: out <= 12'h222;
      20'h06178: out <= 12'h000;
      20'h06179: out <= 12'h000;
      20'h0617a: out <= 12'h000;
      20'h0617b: out <= 12'h666;
      20'h0617c: out <= 12'h666;
      20'h0617d: out <= 12'hbbb;
      20'h0617e: out <= 12'hfff;
      20'h0617f: out <= 12'h666;
      20'h06180: out <= 12'hbbb;
      20'h06181: out <= 12'hfff;
      20'h06182: out <= 12'h666;
      20'h06183: out <= 12'hbbb;
      20'h06184: out <= 12'h666;
      20'h06185: out <= 12'hbbb;
      20'h06186: out <= 12'h000;
      20'h06187: out <= 12'h000;
      20'h06188: out <= 12'h222;
      20'h06189: out <= 12'h222;
      20'h0618a: out <= 12'h222;
      20'h0618b: out <= 12'hbbb;
      20'h0618c: out <= 12'h666;
      20'h0618d: out <= 12'hbbb;
      20'h0618e: out <= 12'hfff;
      20'h0618f: out <= 12'h666;
      20'h06190: out <= 12'hbbb;
      20'h06191: out <= 12'hfff;
      20'h06192: out <= 12'h666;
      20'h06193: out <= 12'hbbb;
      20'h06194: out <= 12'h666;
      20'h06195: out <= 12'h666;
      20'h06196: out <= 12'h222;
      20'h06197: out <= 12'h222;
      20'h06198: out <= 12'h000;
      20'h06199: out <= 12'h000;
      20'h0619a: out <= 12'h000;
      20'h0619b: out <= 12'h666;
      20'h0619c: out <= 12'hbbb;
      20'h0619d: out <= 12'h666;
      20'h0619e: out <= 12'hfff;
      20'h0619f: out <= 12'h666;
      20'h061a0: out <= 12'h666;
      20'h061a1: out <= 12'h666;
      20'h061a2: out <= 12'h666;
      20'h061a3: out <= 12'h666;
      20'h061a4: out <= 12'h666;
      20'h061a5: out <= 12'hbbb;
      20'h061a6: out <= 12'h666;
      20'h061a7: out <= 12'h000;
      20'h061a8: out <= 12'h222;
      20'h061a9: out <= 12'h222;
      20'h061aa: out <= 12'h222;
      20'h061ab: out <= 12'h666;
      20'h061ac: out <= 12'hbbb;
      20'h061ad: out <= 12'h666;
      20'h061ae: out <= 12'hfff;
      20'h061af: out <= 12'h666;
      20'h061b0: out <= 12'h666;
      20'h061b1: out <= 12'h666;
      20'h061b2: out <= 12'h666;
      20'h061b3: out <= 12'h666;
      20'h061b4: out <= 12'h666;
      20'h061b5: out <= 12'hbbb;
      20'h061b6: out <= 12'h666;
      20'h061b7: out <= 12'h222;
      20'h061b8: out <= 12'h000;
      20'h061b9: out <= 12'h000;
      20'h061ba: out <= 12'h000;
      20'h061bb: out <= 12'hbbb;
      20'h061bc: out <= 12'h666;
      20'h061bd: out <= 12'h666;
      20'h061be: out <= 12'hfff;
      20'h061bf: out <= 12'hfff;
      20'h061c0: out <= 12'hfff;
      20'h061c1: out <= 12'hfff;
      20'h061c2: out <= 12'hfff;
      20'h061c3: out <= 12'h666;
      20'h061c4: out <= 12'h666;
      20'h061c5: out <= 12'h666;
      20'h061c6: out <= 12'h000;
      20'h061c7: out <= 12'h000;
      20'h061c8: out <= 12'h222;
      20'h061c9: out <= 12'h222;
      20'h061ca: out <= 12'h222;
      20'h061cb: out <= 12'h666;
      20'h061cc: out <= 12'h666;
      20'h061cd: out <= 12'h666;
      20'h061ce: out <= 12'hfff;
      20'h061cf: out <= 12'hfff;
      20'h061d0: out <= 12'hfff;
      20'h061d1: out <= 12'hfff;
      20'h061d2: out <= 12'hfff;
      20'h061d3: out <= 12'h666;
      20'h061d4: out <= 12'h666;
      20'h061d5: out <= 12'hbbb;
      20'h061d6: out <= 12'h222;
      20'h061d7: out <= 12'h222;
      20'h061d8: out <= 12'h603;
      20'h061d9: out <= 12'h603;
      20'h061da: out <= 12'h603;
      20'h061db: out <= 12'h603;
      20'h061dc: out <= 12'h603;
      20'h061dd: out <= 12'h603;
      20'h061de: out <= 12'h603;
      20'h061df: out <= 12'h603;
      20'h061e0: out <= 12'h603;
      20'h061e1: out <= 12'h603;
      20'h061e2: out <= 12'h603;
      20'h061e3: out <= 12'h603;
      20'h061e4: out <= 12'h603;
      20'h061e5: out <= 12'h603;
      20'h061e6: out <= 12'h603;
      20'h061e7: out <= 12'h603;
      20'h061e8: out <= 12'h603;
      20'h061e9: out <= 12'h603;
      20'h061ea: out <= 12'h603;
      20'h061eb: out <= 12'h603;
      20'h061ec: out <= 12'h603;
      20'h061ed: out <= 12'h603;
      20'h061ee: out <= 12'h603;
      20'h061ef: out <= 12'h603;
      20'h061f0: out <= 12'h603;
      20'h061f1: out <= 12'h603;
      20'h061f2: out <= 12'h603;
      20'h061f3: out <= 12'h603;
      20'h061f4: out <= 12'h603;
      20'h061f5: out <= 12'h603;
      20'h061f6: out <= 12'h603;
      20'h061f7: out <= 12'h603;
      20'h061f8: out <= 12'h603;
      20'h061f9: out <= 12'h603;
      20'h061fa: out <= 12'h603;
      20'h061fb: out <= 12'h603;
      20'h061fc: out <= 12'h603;
      20'h061fd: out <= 12'h603;
      20'h061fe: out <= 12'h603;
      20'h061ff: out <= 12'h603;
      20'h06200: out <= 12'h603;
      20'h06201: out <= 12'h603;
      20'h06202: out <= 12'h603;
      20'h06203: out <= 12'h603;
      20'h06204: out <= 12'h603;
      20'h06205: out <= 12'h603;
      20'h06206: out <= 12'h603;
      20'h06207: out <= 12'h603;
      20'h06208: out <= 12'h603;
      20'h06209: out <= 12'h603;
      20'h0620a: out <= 12'h603;
      20'h0620b: out <= 12'h603;
      20'h0620c: out <= 12'h603;
      20'h0620d: out <= 12'h603;
      20'h0620e: out <= 12'h603;
      20'h0620f: out <= 12'h603;
      20'h06210: out <= 12'h603;
      20'h06211: out <= 12'h603;
      20'h06212: out <= 12'h603;
      20'h06213: out <= 12'h603;
      20'h06214: out <= 12'h603;
      20'h06215: out <= 12'h603;
      20'h06216: out <= 12'h603;
      20'h06217: out <= 12'h603;
      20'h06218: out <= 12'h603;
      20'h06219: out <= 12'h603;
      20'h0621a: out <= 12'h603;
      20'h0621b: out <= 12'h603;
      20'h0621c: out <= 12'h603;
      20'h0621d: out <= 12'h603;
      20'h0621e: out <= 12'h603;
      20'h0621f: out <= 12'h603;
      20'h06220: out <= 12'h603;
      20'h06221: out <= 12'h603;
      20'h06222: out <= 12'h603;
      20'h06223: out <= 12'h603;
      20'h06224: out <= 12'h603;
      20'h06225: out <= 12'h603;
      20'h06226: out <= 12'h603;
      20'h06227: out <= 12'h603;
      20'h06228: out <= 12'h603;
      20'h06229: out <= 12'h603;
      20'h0622a: out <= 12'h603;
      20'h0622b: out <= 12'h603;
      20'h0622c: out <= 12'h603;
      20'h0622d: out <= 12'h603;
      20'h0622e: out <= 12'h603;
      20'h0622f: out <= 12'h603;
      20'h06230: out <= 12'hee9;
      20'h06231: out <= 12'hf87;
      20'h06232: out <= 12'hf87;
      20'h06233: out <= 12'hf87;
      20'h06234: out <= 12'hf87;
      20'h06235: out <= 12'hf87;
      20'h06236: out <= 12'hf87;
      20'h06237: out <= 12'hb27;
      20'h06238: out <= 12'h000;
      20'h06239: out <= 12'h000;
      20'h0623a: out <= 12'h000;
      20'h0623b: out <= 12'h000;
      20'h0623c: out <= 12'h000;
      20'h0623d: out <= 12'h000;
      20'h0623e: out <= 12'h000;
      20'h0623f: out <= 12'h000;
      20'h06240: out <= 12'hfa9;
      20'h06241: out <= 12'hfa9;
      20'h06242: out <= 12'hfa9;
      20'h06243: out <= 12'hfa9;
      20'h06244: out <= 12'hfa9;
      20'h06245: out <= 12'hfa9;
      20'h06246: out <= 12'hfa9;
      20'h06247: out <= 12'hfa9;
      20'h06248: out <= 12'hf76;
      20'h06249: out <= 12'hf76;
      20'h0624a: out <= 12'hf76;
      20'h0624b: out <= 12'hf76;
      20'h0624c: out <= 12'hf76;
      20'h0624d: out <= 12'hf76;
      20'h0624e: out <= 12'hf76;
      20'h0624f: out <= 12'hf76;
      20'h06250: out <= 12'hfa9;
      20'h06251: out <= 12'hfa9;
      20'h06252: out <= 12'hfa9;
      20'h06253: out <= 12'hfa9;
      20'h06254: out <= 12'hfa9;
      20'h06255: out <= 12'hfa9;
      20'h06256: out <= 12'hfa9;
      20'h06257: out <= 12'hfa9;
      20'h06258: out <= 12'hf76;
      20'h06259: out <= 12'hf76;
      20'h0625a: out <= 12'hf76;
      20'h0625b: out <= 12'hf76;
      20'h0625c: out <= 12'hf76;
      20'h0625d: out <= 12'hf76;
      20'h0625e: out <= 12'hf76;
      20'h0625f: out <= 12'hf76;
      20'h06260: out <= 12'hfa9;
      20'h06261: out <= 12'hfa9;
      20'h06262: out <= 12'hfa9;
      20'h06263: out <= 12'hfa9;
      20'h06264: out <= 12'hfa9;
      20'h06265: out <= 12'hfa9;
      20'h06266: out <= 12'hfa9;
      20'h06267: out <= 12'hfa9;
      20'h06268: out <= 12'h000;
      20'h06269: out <= 12'h000;
      20'h0626a: out <= 12'h000;
      20'h0626b: out <= 12'h000;
      20'h0626c: out <= 12'h000;
      20'h0626d: out <= 12'h000;
      20'h0626e: out <= 12'h000;
      20'h0626f: out <= 12'h000;
      20'h06270: out <= 12'h000;
      20'h06271: out <= 12'h000;
      20'h06272: out <= 12'h666;
      20'h06273: out <= 12'hbbb;
      20'h06274: out <= 12'hbbb;
      20'h06275: out <= 12'hbbb;
      20'h06276: out <= 12'hbbb;
      20'h06277: out <= 12'hbbb;
      20'h06278: out <= 12'hbbb;
      20'h06279: out <= 12'h666;
      20'h0627a: out <= 12'hbbb;
      20'h0627b: out <= 12'hfff;
      20'h0627c: out <= 12'h666;
      20'h0627d: out <= 12'h000;
      20'h0627e: out <= 12'h000;
      20'h0627f: out <= 12'h000;
      20'h06280: out <= 12'h222;
      20'h06281: out <= 12'h222;
      20'h06282: out <= 12'h666;
      20'h06283: out <= 12'hbbb;
      20'h06284: out <= 12'hbbb;
      20'h06285: out <= 12'hbbb;
      20'h06286: out <= 12'hbbb;
      20'h06287: out <= 12'hbbb;
      20'h06288: out <= 12'hbbb;
      20'h06289: out <= 12'h666;
      20'h0628a: out <= 12'hbbb;
      20'h0628b: out <= 12'hfff;
      20'h0628c: out <= 12'h666;
      20'h0628d: out <= 12'h222;
      20'h0628e: out <= 12'h222;
      20'h0628f: out <= 12'h222;
      20'h06290: out <= 12'h000;
      20'h06291: out <= 12'h000;
      20'h06292: out <= 12'h000;
      20'h06293: out <= 12'hbbb;
      20'h06294: out <= 12'h666;
      20'h06295: out <= 12'hbbb;
      20'h06296: out <= 12'hfff;
      20'h06297: out <= 12'h666;
      20'h06298: out <= 12'hfff;
      20'h06299: out <= 12'hfff;
      20'h0629a: out <= 12'h666;
      20'h0629b: out <= 12'hbbb;
      20'h0629c: out <= 12'h666;
      20'h0629d: out <= 12'h666;
      20'h0629e: out <= 12'h000;
      20'h0629f: out <= 12'h000;
      20'h062a0: out <= 12'h222;
      20'h062a1: out <= 12'h222;
      20'h062a2: out <= 12'h222;
      20'h062a3: out <= 12'h666;
      20'h062a4: out <= 12'h666;
      20'h062a5: out <= 12'hbbb;
      20'h062a6: out <= 12'hfff;
      20'h062a7: out <= 12'h666;
      20'h062a8: out <= 12'hfff;
      20'h062a9: out <= 12'hfff;
      20'h062aa: out <= 12'h666;
      20'h062ab: out <= 12'hbbb;
      20'h062ac: out <= 12'h666;
      20'h062ad: out <= 12'hbbb;
      20'h062ae: out <= 12'h222;
      20'h062af: out <= 12'h222;
      20'h062b0: out <= 12'h000;
      20'h062b1: out <= 12'h000;
      20'h062b2: out <= 12'h000;
      20'h062b3: out <= 12'h666;
      20'h062b4: out <= 12'hfff;
      20'h062b5: out <= 12'hbbb;
      20'h062b6: out <= 12'h666;
      20'h062b7: out <= 12'hbbb;
      20'h062b8: out <= 12'hbbb;
      20'h062b9: out <= 12'hbbb;
      20'h062ba: out <= 12'hbbb;
      20'h062bb: out <= 12'hbbb;
      20'h062bc: out <= 12'hbbb;
      20'h062bd: out <= 12'h666;
      20'h062be: out <= 12'h000;
      20'h062bf: out <= 12'h000;
      20'h062c0: out <= 12'h222;
      20'h062c1: out <= 12'h222;
      20'h062c2: out <= 12'h222;
      20'h062c3: out <= 12'h666;
      20'h062c4: out <= 12'hfff;
      20'h062c5: out <= 12'hbbb;
      20'h062c6: out <= 12'h666;
      20'h062c7: out <= 12'hbbb;
      20'h062c8: out <= 12'hbbb;
      20'h062c9: out <= 12'hbbb;
      20'h062ca: out <= 12'hbbb;
      20'h062cb: out <= 12'hbbb;
      20'h062cc: out <= 12'hbbb;
      20'h062cd: out <= 12'h666;
      20'h062ce: out <= 12'h222;
      20'h062cf: out <= 12'h222;
      20'h062d0: out <= 12'h000;
      20'h062d1: out <= 12'h000;
      20'h062d2: out <= 12'h000;
      20'h062d3: out <= 12'h666;
      20'h062d4: out <= 12'h666;
      20'h062d5: out <= 12'hbbb;
      20'h062d6: out <= 12'h666;
      20'h062d7: out <= 12'h666;
      20'h062d8: out <= 12'hbbb;
      20'h062d9: out <= 12'h666;
      20'h062da: out <= 12'h666;
      20'h062db: out <= 12'hbbb;
      20'h062dc: out <= 12'h666;
      20'h062dd: out <= 12'hbbb;
      20'h062de: out <= 12'h000;
      20'h062df: out <= 12'h000;
      20'h062e0: out <= 12'h222;
      20'h062e1: out <= 12'h222;
      20'h062e2: out <= 12'h222;
      20'h062e3: out <= 12'hbbb;
      20'h062e4: out <= 12'h666;
      20'h062e5: out <= 12'hbbb;
      20'h062e6: out <= 12'h666;
      20'h062e7: out <= 12'h666;
      20'h062e8: out <= 12'hbbb;
      20'h062e9: out <= 12'h666;
      20'h062ea: out <= 12'h666;
      20'h062eb: out <= 12'hbbb;
      20'h062ec: out <= 12'h666;
      20'h062ed: out <= 12'h666;
      20'h062ee: out <= 12'h222;
      20'h062ef: out <= 12'h222;
      20'h062f0: out <= 12'h603;
      20'h062f1: out <= 12'h603;
      20'h062f2: out <= 12'h603;
      20'h062f3: out <= 12'h603;
      20'h062f4: out <= 12'h603;
      20'h062f5: out <= 12'h603;
      20'h062f6: out <= 12'h603;
      20'h062f7: out <= 12'h603;
      20'h062f8: out <= 12'h603;
      20'h062f9: out <= 12'h603;
      20'h062fa: out <= 12'h603;
      20'h062fb: out <= 12'h603;
      20'h062fc: out <= 12'h603;
      20'h062fd: out <= 12'h603;
      20'h062fe: out <= 12'h603;
      20'h062ff: out <= 12'h603;
      20'h06300: out <= 12'h603;
      20'h06301: out <= 12'h603;
      20'h06302: out <= 12'h603;
      20'h06303: out <= 12'h603;
      20'h06304: out <= 12'h603;
      20'h06305: out <= 12'h603;
      20'h06306: out <= 12'h603;
      20'h06307: out <= 12'h603;
      20'h06308: out <= 12'h603;
      20'h06309: out <= 12'h603;
      20'h0630a: out <= 12'h603;
      20'h0630b: out <= 12'h603;
      20'h0630c: out <= 12'h603;
      20'h0630d: out <= 12'h603;
      20'h0630e: out <= 12'h603;
      20'h0630f: out <= 12'h603;
      20'h06310: out <= 12'h603;
      20'h06311: out <= 12'h603;
      20'h06312: out <= 12'h603;
      20'h06313: out <= 12'h603;
      20'h06314: out <= 12'h603;
      20'h06315: out <= 12'h603;
      20'h06316: out <= 12'h603;
      20'h06317: out <= 12'h603;
      20'h06318: out <= 12'h603;
      20'h06319: out <= 12'h603;
      20'h0631a: out <= 12'h603;
      20'h0631b: out <= 12'h603;
      20'h0631c: out <= 12'h603;
      20'h0631d: out <= 12'h603;
      20'h0631e: out <= 12'h603;
      20'h0631f: out <= 12'h603;
      20'h06320: out <= 12'h603;
      20'h06321: out <= 12'h603;
      20'h06322: out <= 12'h603;
      20'h06323: out <= 12'h603;
      20'h06324: out <= 12'h603;
      20'h06325: out <= 12'h603;
      20'h06326: out <= 12'h603;
      20'h06327: out <= 12'h603;
      20'h06328: out <= 12'h603;
      20'h06329: out <= 12'h603;
      20'h0632a: out <= 12'h603;
      20'h0632b: out <= 12'h603;
      20'h0632c: out <= 12'h603;
      20'h0632d: out <= 12'h603;
      20'h0632e: out <= 12'h603;
      20'h0632f: out <= 12'h603;
      20'h06330: out <= 12'h603;
      20'h06331: out <= 12'h603;
      20'h06332: out <= 12'h603;
      20'h06333: out <= 12'h603;
      20'h06334: out <= 12'h603;
      20'h06335: out <= 12'h603;
      20'h06336: out <= 12'h603;
      20'h06337: out <= 12'h603;
      20'h06338: out <= 12'h603;
      20'h06339: out <= 12'h603;
      20'h0633a: out <= 12'h603;
      20'h0633b: out <= 12'h603;
      20'h0633c: out <= 12'h603;
      20'h0633d: out <= 12'h603;
      20'h0633e: out <= 12'h603;
      20'h0633f: out <= 12'h603;
      20'h06340: out <= 12'h603;
      20'h06341: out <= 12'h603;
      20'h06342: out <= 12'h603;
      20'h06343: out <= 12'h603;
      20'h06344: out <= 12'h603;
      20'h06345: out <= 12'h603;
      20'h06346: out <= 12'h603;
      20'h06347: out <= 12'h603;
      20'h06348: out <= 12'hee9;
      20'h06349: out <= 12'hf87;
      20'h0634a: out <= 12'hee9;
      20'h0634b: out <= 12'hee9;
      20'h0634c: out <= 12'hee9;
      20'h0634d: out <= 12'hb27;
      20'h0634e: out <= 12'hf87;
      20'h0634f: out <= 12'hb27;
      20'h06350: out <= 12'h000;
      20'h06351: out <= 12'h000;
      20'h06352: out <= 12'h000;
      20'h06353: out <= 12'h000;
      20'h06354: out <= 12'h000;
      20'h06355: out <= 12'h000;
      20'h06356: out <= 12'h000;
      20'h06357: out <= 12'h000;
      20'h06358: out <= 12'hfa9;
      20'h06359: out <= 12'hfa9;
      20'h0635a: out <= 12'hfa9;
      20'h0635b: out <= 12'hfa9;
      20'h0635c: out <= 12'hfa9;
      20'h0635d: out <= 12'hfa9;
      20'h0635e: out <= 12'hfa9;
      20'h0635f: out <= 12'hfa9;
      20'h06360: out <= 12'hf76;
      20'h06361: out <= 12'hf76;
      20'h06362: out <= 12'hf76;
      20'h06363: out <= 12'hf76;
      20'h06364: out <= 12'hf76;
      20'h06365: out <= 12'hf76;
      20'h06366: out <= 12'hf76;
      20'h06367: out <= 12'hf76;
      20'h06368: out <= 12'hfa9;
      20'h06369: out <= 12'hfa9;
      20'h0636a: out <= 12'hfa9;
      20'h0636b: out <= 12'hfa9;
      20'h0636c: out <= 12'hfa9;
      20'h0636d: out <= 12'hfa9;
      20'h0636e: out <= 12'hfa9;
      20'h0636f: out <= 12'hfa9;
      20'h06370: out <= 12'hf76;
      20'h06371: out <= 12'hf76;
      20'h06372: out <= 12'hf76;
      20'h06373: out <= 12'hf76;
      20'h06374: out <= 12'hf76;
      20'h06375: out <= 12'hf76;
      20'h06376: out <= 12'hf76;
      20'h06377: out <= 12'hf76;
      20'h06378: out <= 12'hfa9;
      20'h06379: out <= 12'hfa9;
      20'h0637a: out <= 12'hfa9;
      20'h0637b: out <= 12'hfa9;
      20'h0637c: out <= 12'hfa9;
      20'h0637d: out <= 12'hfa9;
      20'h0637e: out <= 12'hfa9;
      20'h0637f: out <= 12'hfa9;
      20'h06380: out <= 12'h000;
      20'h06381: out <= 12'h000;
      20'h06382: out <= 12'h000;
      20'h06383: out <= 12'h000;
      20'h06384: out <= 12'h000;
      20'h06385: out <= 12'h000;
      20'h06386: out <= 12'h000;
      20'h06387: out <= 12'h000;
      20'h06388: out <= 12'h000;
      20'h06389: out <= 12'h000;
      20'h0638a: out <= 12'h000;
      20'h0638b: out <= 12'h666;
      20'h0638c: out <= 12'h666;
      20'h0638d: out <= 12'h666;
      20'h0638e: out <= 12'h666;
      20'h0638f: out <= 12'h666;
      20'h06390: out <= 12'h666;
      20'h06391: out <= 12'h666;
      20'h06392: out <= 12'h666;
      20'h06393: out <= 12'h666;
      20'h06394: out <= 12'h000;
      20'h06395: out <= 12'h000;
      20'h06396: out <= 12'h000;
      20'h06397: out <= 12'h000;
      20'h06398: out <= 12'h222;
      20'h06399: out <= 12'h222;
      20'h0639a: out <= 12'h222;
      20'h0639b: out <= 12'h666;
      20'h0639c: out <= 12'h666;
      20'h0639d: out <= 12'h666;
      20'h0639e: out <= 12'h666;
      20'h0639f: out <= 12'h666;
      20'h063a0: out <= 12'h666;
      20'h063a1: out <= 12'h666;
      20'h063a2: out <= 12'h666;
      20'h063a3: out <= 12'h666;
      20'h063a4: out <= 12'h222;
      20'h063a5: out <= 12'h222;
      20'h063a6: out <= 12'h222;
      20'h063a7: out <= 12'h222;
      20'h063a8: out <= 12'h000;
      20'h063a9: out <= 12'h000;
      20'h063aa: out <= 12'h000;
      20'h063ab: out <= 12'h666;
      20'h063ac: out <= 12'h666;
      20'h063ad: out <= 12'hbbb;
      20'h063ae: out <= 12'hfff;
      20'h063af: out <= 12'hbbb;
      20'h063b0: out <= 12'hbbb;
      20'h063b1: out <= 12'hbbb;
      20'h063b2: out <= 12'h666;
      20'h063b3: out <= 12'hbbb;
      20'h063b4: out <= 12'h666;
      20'h063b5: out <= 12'hbbb;
      20'h063b6: out <= 12'h000;
      20'h063b7: out <= 12'h000;
      20'h063b8: out <= 12'h222;
      20'h063b9: out <= 12'h222;
      20'h063ba: out <= 12'h222;
      20'h063bb: out <= 12'hbbb;
      20'h063bc: out <= 12'h666;
      20'h063bd: out <= 12'hbbb;
      20'h063be: out <= 12'hfff;
      20'h063bf: out <= 12'hbbb;
      20'h063c0: out <= 12'hbbb;
      20'h063c1: out <= 12'hbbb;
      20'h063c2: out <= 12'h666;
      20'h063c3: out <= 12'hbbb;
      20'h063c4: out <= 12'h666;
      20'h063c5: out <= 12'h666;
      20'h063c6: out <= 12'h222;
      20'h063c7: out <= 12'h222;
      20'h063c8: out <= 12'h000;
      20'h063c9: out <= 12'h000;
      20'h063ca: out <= 12'h000;
      20'h063cb: out <= 12'h000;
      20'h063cc: out <= 12'h666;
      20'h063cd: out <= 12'h666;
      20'h063ce: out <= 12'h666;
      20'h063cf: out <= 12'h666;
      20'h063d0: out <= 12'h666;
      20'h063d1: out <= 12'h666;
      20'h063d2: out <= 12'h666;
      20'h063d3: out <= 12'h666;
      20'h063d4: out <= 12'h666;
      20'h063d5: out <= 12'h000;
      20'h063d6: out <= 12'h000;
      20'h063d7: out <= 12'h000;
      20'h063d8: out <= 12'h222;
      20'h063d9: out <= 12'h222;
      20'h063da: out <= 12'h222;
      20'h063db: out <= 12'h222;
      20'h063dc: out <= 12'h666;
      20'h063dd: out <= 12'h666;
      20'h063de: out <= 12'h666;
      20'h063df: out <= 12'h666;
      20'h063e0: out <= 12'h666;
      20'h063e1: out <= 12'h666;
      20'h063e2: out <= 12'h666;
      20'h063e3: out <= 12'h666;
      20'h063e4: out <= 12'h666;
      20'h063e5: out <= 12'h222;
      20'h063e6: out <= 12'h222;
      20'h063e7: out <= 12'h222;
      20'h063e8: out <= 12'h000;
      20'h063e9: out <= 12'h000;
      20'h063ea: out <= 12'h000;
      20'h063eb: out <= 12'hfff;
      20'h063ec: out <= 12'h666;
      20'h063ed: out <= 12'hfff;
      20'h063ee: out <= 12'hbbb;
      20'h063ef: out <= 12'h666;
      20'h063f0: out <= 12'hbbb;
      20'h063f1: out <= 12'h666;
      20'h063f2: out <= 12'hbbb;
      20'h063f3: out <= 12'hfff;
      20'h063f4: out <= 12'h666;
      20'h063f5: out <= 12'hfff;
      20'h063f6: out <= 12'h000;
      20'h063f7: out <= 12'h000;
      20'h063f8: out <= 12'h222;
      20'h063f9: out <= 12'h222;
      20'h063fa: out <= 12'h222;
      20'h063fb: out <= 12'hfff;
      20'h063fc: out <= 12'h666;
      20'h063fd: out <= 12'hfff;
      20'h063fe: out <= 12'hbbb;
      20'h063ff: out <= 12'h666;
      20'h06400: out <= 12'hbbb;
      20'h06401: out <= 12'h666;
      20'h06402: out <= 12'hbbb;
      20'h06403: out <= 12'hfff;
      20'h06404: out <= 12'h666;
      20'h06405: out <= 12'hfff;
      20'h06406: out <= 12'h222;
      20'h06407: out <= 12'h222;
      20'h06408: out <= 12'h603;
      20'h06409: out <= 12'h603;
      20'h0640a: out <= 12'h603;
      20'h0640b: out <= 12'h603;
      20'h0640c: out <= 12'h603;
      20'h0640d: out <= 12'h603;
      20'h0640e: out <= 12'h603;
      20'h0640f: out <= 12'h603;
      20'h06410: out <= 12'h603;
      20'h06411: out <= 12'h603;
      20'h06412: out <= 12'h603;
      20'h06413: out <= 12'h603;
      20'h06414: out <= 12'h603;
      20'h06415: out <= 12'h603;
      20'h06416: out <= 12'h603;
      20'h06417: out <= 12'h603;
      20'h06418: out <= 12'h603;
      20'h06419: out <= 12'h603;
      20'h0641a: out <= 12'h603;
      20'h0641b: out <= 12'h603;
      20'h0641c: out <= 12'h603;
      20'h0641d: out <= 12'h603;
      20'h0641e: out <= 12'h603;
      20'h0641f: out <= 12'h603;
      20'h06420: out <= 12'h603;
      20'h06421: out <= 12'h603;
      20'h06422: out <= 12'h603;
      20'h06423: out <= 12'h603;
      20'h06424: out <= 12'h603;
      20'h06425: out <= 12'h603;
      20'h06426: out <= 12'h603;
      20'h06427: out <= 12'h603;
      20'h06428: out <= 12'h603;
      20'h06429: out <= 12'h603;
      20'h0642a: out <= 12'h603;
      20'h0642b: out <= 12'h603;
      20'h0642c: out <= 12'h603;
      20'h0642d: out <= 12'h603;
      20'h0642e: out <= 12'h603;
      20'h0642f: out <= 12'h603;
      20'h06430: out <= 12'h603;
      20'h06431: out <= 12'h603;
      20'h06432: out <= 12'h603;
      20'h06433: out <= 12'h603;
      20'h06434: out <= 12'h603;
      20'h06435: out <= 12'h603;
      20'h06436: out <= 12'h603;
      20'h06437: out <= 12'h603;
      20'h06438: out <= 12'h603;
      20'h06439: out <= 12'h603;
      20'h0643a: out <= 12'h603;
      20'h0643b: out <= 12'h603;
      20'h0643c: out <= 12'h603;
      20'h0643d: out <= 12'h603;
      20'h0643e: out <= 12'h603;
      20'h0643f: out <= 12'h603;
      20'h06440: out <= 12'h603;
      20'h06441: out <= 12'h603;
      20'h06442: out <= 12'h603;
      20'h06443: out <= 12'h603;
      20'h06444: out <= 12'h603;
      20'h06445: out <= 12'h603;
      20'h06446: out <= 12'h603;
      20'h06447: out <= 12'h603;
      20'h06448: out <= 12'h603;
      20'h06449: out <= 12'h603;
      20'h0644a: out <= 12'h603;
      20'h0644b: out <= 12'h603;
      20'h0644c: out <= 12'h603;
      20'h0644d: out <= 12'h603;
      20'h0644e: out <= 12'h603;
      20'h0644f: out <= 12'h603;
      20'h06450: out <= 12'h603;
      20'h06451: out <= 12'h603;
      20'h06452: out <= 12'h603;
      20'h06453: out <= 12'h603;
      20'h06454: out <= 12'h603;
      20'h06455: out <= 12'h603;
      20'h06456: out <= 12'h603;
      20'h06457: out <= 12'h603;
      20'h06458: out <= 12'h603;
      20'h06459: out <= 12'h603;
      20'h0645a: out <= 12'h603;
      20'h0645b: out <= 12'h603;
      20'h0645c: out <= 12'h603;
      20'h0645d: out <= 12'h603;
      20'h0645e: out <= 12'h603;
      20'h0645f: out <= 12'h603;
      20'h06460: out <= 12'hee9;
      20'h06461: out <= 12'hf87;
      20'h06462: out <= 12'hee9;
      20'h06463: out <= 12'hf87;
      20'h06464: out <= 12'hf87;
      20'h06465: out <= 12'hb27;
      20'h06466: out <= 12'hf87;
      20'h06467: out <= 12'hb27;
      20'h06468: out <= 12'h000;
      20'h06469: out <= 12'h000;
      20'h0646a: out <= 12'h000;
      20'h0646b: out <= 12'h000;
      20'h0646c: out <= 12'h000;
      20'h0646d: out <= 12'h000;
      20'h0646e: out <= 12'h000;
      20'h0646f: out <= 12'h000;
      20'h06470: out <= 12'hfa9;
      20'h06471: out <= 12'hfa9;
      20'h06472: out <= 12'hfa9;
      20'h06473: out <= 12'hfa9;
      20'h06474: out <= 12'hfa9;
      20'h06475: out <= 12'hfa9;
      20'h06476: out <= 12'hfa9;
      20'h06477: out <= 12'hfa9;
      20'h06478: out <= 12'hf76;
      20'h06479: out <= 12'hf76;
      20'h0647a: out <= 12'hf76;
      20'h0647b: out <= 12'hf76;
      20'h0647c: out <= 12'hf76;
      20'h0647d: out <= 12'hf76;
      20'h0647e: out <= 12'hf76;
      20'h0647f: out <= 12'hf76;
      20'h06480: out <= 12'hfa9;
      20'h06481: out <= 12'hfa9;
      20'h06482: out <= 12'hfa9;
      20'h06483: out <= 12'hfa9;
      20'h06484: out <= 12'hfa9;
      20'h06485: out <= 12'hfa9;
      20'h06486: out <= 12'hfa9;
      20'h06487: out <= 12'hfa9;
      20'h06488: out <= 12'hf76;
      20'h06489: out <= 12'hf76;
      20'h0648a: out <= 12'hf76;
      20'h0648b: out <= 12'hf76;
      20'h0648c: out <= 12'hf76;
      20'h0648d: out <= 12'hf76;
      20'h0648e: out <= 12'hf76;
      20'h0648f: out <= 12'hf76;
      20'h06490: out <= 12'hfa9;
      20'h06491: out <= 12'hfa9;
      20'h06492: out <= 12'hfa9;
      20'h06493: out <= 12'hfa9;
      20'h06494: out <= 12'hfa9;
      20'h06495: out <= 12'hfa9;
      20'h06496: out <= 12'hfa9;
      20'h06497: out <= 12'hfa9;
      20'h06498: out <= 12'h000;
      20'h06499: out <= 12'h000;
      20'h0649a: out <= 12'h000;
      20'h0649b: out <= 12'h000;
      20'h0649c: out <= 12'h000;
      20'h0649d: out <= 12'h000;
      20'h0649e: out <= 12'h000;
      20'h0649f: out <= 12'h000;
      20'h064a0: out <= 12'h000;
      20'h064a1: out <= 12'h000;
      20'h064a2: out <= 12'h000;
      20'h064a3: out <= 12'hfff;
      20'h064a4: out <= 12'hbbb;
      20'h064a5: out <= 12'h666;
      20'h064a6: out <= 12'hbbb;
      20'h064a7: out <= 12'h666;
      20'h064a8: out <= 12'hbbb;
      20'h064a9: out <= 12'h666;
      20'h064aa: out <= 12'hbbb;
      20'h064ab: out <= 12'hfff;
      20'h064ac: out <= 12'h000;
      20'h064ad: out <= 12'h000;
      20'h064ae: out <= 12'h000;
      20'h064af: out <= 12'h000;
      20'h064b0: out <= 12'h222;
      20'h064b1: out <= 12'h222;
      20'h064b2: out <= 12'h222;
      20'h064b3: out <= 12'hfff;
      20'h064b4: out <= 12'h666;
      20'h064b5: out <= 12'hbbb;
      20'h064b6: out <= 12'h666;
      20'h064b7: out <= 12'hbbb;
      20'h064b8: out <= 12'h666;
      20'h064b9: out <= 12'hbbb;
      20'h064ba: out <= 12'h666;
      20'h064bb: out <= 12'hfff;
      20'h064bc: out <= 12'h222;
      20'h064bd: out <= 12'h222;
      20'h064be: out <= 12'h222;
      20'h064bf: out <= 12'h222;
      20'h064c0: out <= 12'h000;
      20'h064c1: out <= 12'h000;
      20'h064c2: out <= 12'h000;
      20'h064c3: out <= 12'hfff;
      20'h064c4: out <= 12'h666;
      20'h064c5: out <= 12'hbbb;
      20'h064c6: out <= 12'hfff;
      20'h064c7: out <= 12'h666;
      20'h064c8: out <= 12'h666;
      20'h064c9: out <= 12'h666;
      20'h064ca: out <= 12'h666;
      20'h064cb: out <= 12'hbbb;
      20'h064cc: out <= 12'h666;
      20'h064cd: out <= 12'hfff;
      20'h064ce: out <= 12'h000;
      20'h064cf: out <= 12'h000;
      20'h064d0: out <= 12'h222;
      20'h064d1: out <= 12'h222;
      20'h064d2: out <= 12'h222;
      20'h064d3: out <= 12'hfff;
      20'h064d4: out <= 12'h666;
      20'h064d5: out <= 12'hbbb;
      20'h064d6: out <= 12'hfff;
      20'h064d7: out <= 12'h666;
      20'h064d8: out <= 12'h666;
      20'h064d9: out <= 12'h666;
      20'h064da: out <= 12'h666;
      20'h064db: out <= 12'hbbb;
      20'h064dc: out <= 12'h666;
      20'h064dd: out <= 12'hfff;
      20'h064de: out <= 12'h222;
      20'h064df: out <= 12'h222;
      20'h064e0: out <= 12'h000;
      20'h064e1: out <= 12'h000;
      20'h064e2: out <= 12'h000;
      20'h064e3: out <= 12'h000;
      20'h064e4: out <= 12'hfff;
      20'h064e5: out <= 12'hbbb;
      20'h064e6: out <= 12'h666;
      20'h064e7: out <= 12'hbbb;
      20'h064e8: out <= 12'h666;
      20'h064e9: out <= 12'hbbb;
      20'h064ea: out <= 12'h666;
      20'h064eb: out <= 12'hbbb;
      20'h064ec: out <= 12'hfff;
      20'h064ed: out <= 12'h000;
      20'h064ee: out <= 12'h000;
      20'h064ef: out <= 12'h000;
      20'h064f0: out <= 12'h222;
      20'h064f1: out <= 12'h222;
      20'h064f2: out <= 12'h222;
      20'h064f3: out <= 12'h222;
      20'h064f4: out <= 12'hfff;
      20'h064f5: out <= 12'h666;
      20'h064f6: out <= 12'hbbb;
      20'h064f7: out <= 12'h666;
      20'h064f8: out <= 12'hbbb;
      20'h064f9: out <= 12'h666;
      20'h064fa: out <= 12'hbbb;
      20'h064fb: out <= 12'h666;
      20'h064fc: out <= 12'hfff;
      20'h064fd: out <= 12'h222;
      20'h064fe: out <= 12'h222;
      20'h064ff: out <= 12'h222;
      20'h06500: out <= 12'h000;
      20'h06501: out <= 12'h000;
      20'h06502: out <= 12'h000;
      20'h06503: out <= 12'h000;
      20'h06504: out <= 12'h000;
      20'h06505: out <= 12'h666;
      20'h06506: out <= 12'h666;
      20'h06507: out <= 12'h666;
      20'h06508: out <= 12'hfff;
      20'h06509: out <= 12'h666;
      20'h0650a: out <= 12'h666;
      20'h0650b: out <= 12'h666;
      20'h0650c: out <= 12'h000;
      20'h0650d: out <= 12'h000;
      20'h0650e: out <= 12'h000;
      20'h0650f: out <= 12'h000;
      20'h06510: out <= 12'h222;
      20'h06511: out <= 12'h222;
      20'h06512: out <= 12'h222;
      20'h06513: out <= 12'h222;
      20'h06514: out <= 12'h222;
      20'h06515: out <= 12'h666;
      20'h06516: out <= 12'h666;
      20'h06517: out <= 12'h666;
      20'h06518: out <= 12'hfff;
      20'h06519: out <= 12'h666;
      20'h0651a: out <= 12'h666;
      20'h0651b: out <= 12'h666;
      20'h0651c: out <= 12'h222;
      20'h0651d: out <= 12'h222;
      20'h0651e: out <= 12'h222;
      20'h0651f: out <= 12'h222;
      20'h06520: out <= 12'h603;
      20'h06521: out <= 12'h603;
      20'h06522: out <= 12'h603;
      20'h06523: out <= 12'h603;
      20'h06524: out <= 12'h603;
      20'h06525: out <= 12'h603;
      20'h06526: out <= 12'h603;
      20'h06527: out <= 12'h603;
      20'h06528: out <= 12'h603;
      20'h06529: out <= 12'h603;
      20'h0652a: out <= 12'h603;
      20'h0652b: out <= 12'h603;
      20'h0652c: out <= 12'h603;
      20'h0652d: out <= 12'h603;
      20'h0652e: out <= 12'h603;
      20'h0652f: out <= 12'h603;
      20'h06530: out <= 12'h603;
      20'h06531: out <= 12'h603;
      20'h06532: out <= 12'h603;
      20'h06533: out <= 12'h603;
      20'h06534: out <= 12'h603;
      20'h06535: out <= 12'h603;
      20'h06536: out <= 12'h603;
      20'h06537: out <= 12'h603;
      20'h06538: out <= 12'h603;
      20'h06539: out <= 12'h603;
      20'h0653a: out <= 12'h603;
      20'h0653b: out <= 12'h603;
      20'h0653c: out <= 12'h603;
      20'h0653d: out <= 12'h603;
      20'h0653e: out <= 12'h603;
      20'h0653f: out <= 12'h603;
      20'h06540: out <= 12'h603;
      20'h06541: out <= 12'h603;
      20'h06542: out <= 12'h603;
      20'h06543: out <= 12'h603;
      20'h06544: out <= 12'h603;
      20'h06545: out <= 12'h603;
      20'h06546: out <= 12'h603;
      20'h06547: out <= 12'h603;
      20'h06548: out <= 12'h603;
      20'h06549: out <= 12'h603;
      20'h0654a: out <= 12'h603;
      20'h0654b: out <= 12'h603;
      20'h0654c: out <= 12'h603;
      20'h0654d: out <= 12'h603;
      20'h0654e: out <= 12'h603;
      20'h0654f: out <= 12'h603;
      20'h06550: out <= 12'h603;
      20'h06551: out <= 12'h603;
      20'h06552: out <= 12'h603;
      20'h06553: out <= 12'h603;
      20'h06554: out <= 12'h603;
      20'h06555: out <= 12'h603;
      20'h06556: out <= 12'h603;
      20'h06557: out <= 12'h603;
      20'h06558: out <= 12'h603;
      20'h06559: out <= 12'h603;
      20'h0655a: out <= 12'h603;
      20'h0655b: out <= 12'h603;
      20'h0655c: out <= 12'h603;
      20'h0655d: out <= 12'h603;
      20'h0655e: out <= 12'h603;
      20'h0655f: out <= 12'h603;
      20'h06560: out <= 12'h603;
      20'h06561: out <= 12'h603;
      20'h06562: out <= 12'h603;
      20'h06563: out <= 12'h603;
      20'h06564: out <= 12'h603;
      20'h06565: out <= 12'h603;
      20'h06566: out <= 12'h603;
      20'h06567: out <= 12'h603;
      20'h06568: out <= 12'h603;
      20'h06569: out <= 12'h603;
      20'h0656a: out <= 12'h603;
      20'h0656b: out <= 12'h603;
      20'h0656c: out <= 12'h603;
      20'h0656d: out <= 12'h603;
      20'h0656e: out <= 12'h603;
      20'h0656f: out <= 12'h603;
      20'h06570: out <= 12'h603;
      20'h06571: out <= 12'h603;
      20'h06572: out <= 12'h603;
      20'h06573: out <= 12'h603;
      20'h06574: out <= 12'h603;
      20'h06575: out <= 12'h603;
      20'h06576: out <= 12'h603;
      20'h06577: out <= 12'h603;
      20'h06578: out <= 12'hee9;
      20'h06579: out <= 12'hf87;
      20'h0657a: out <= 12'hee9;
      20'h0657b: out <= 12'hf87;
      20'h0657c: out <= 12'hf87;
      20'h0657d: out <= 12'hb27;
      20'h0657e: out <= 12'hf87;
      20'h0657f: out <= 12'hb27;
      20'h06580: out <= 12'h000;
      20'h06581: out <= 12'h000;
      20'h06582: out <= 12'h000;
      20'h06583: out <= 12'h000;
      20'h06584: out <= 12'h000;
      20'h06585: out <= 12'h000;
      20'h06586: out <= 12'h000;
      20'h06587: out <= 12'h000;
      20'h06588: out <= 12'hfa9;
      20'h06589: out <= 12'hfa9;
      20'h0658a: out <= 12'hfa9;
      20'h0658b: out <= 12'hfa9;
      20'h0658c: out <= 12'hfa9;
      20'h0658d: out <= 12'hfa9;
      20'h0658e: out <= 12'hfa9;
      20'h0658f: out <= 12'hfa9;
      20'h06590: out <= 12'hf76;
      20'h06591: out <= 12'hf76;
      20'h06592: out <= 12'hf76;
      20'h06593: out <= 12'hf76;
      20'h06594: out <= 12'hf76;
      20'h06595: out <= 12'hf76;
      20'h06596: out <= 12'hf76;
      20'h06597: out <= 12'hf76;
      20'h06598: out <= 12'hfa9;
      20'h06599: out <= 12'hfa9;
      20'h0659a: out <= 12'hfa9;
      20'h0659b: out <= 12'hfa9;
      20'h0659c: out <= 12'hfa9;
      20'h0659d: out <= 12'hfa9;
      20'h0659e: out <= 12'hfa9;
      20'h0659f: out <= 12'hfa9;
      20'h065a0: out <= 12'hf76;
      20'h065a1: out <= 12'hf76;
      20'h065a2: out <= 12'hf76;
      20'h065a3: out <= 12'hf76;
      20'h065a4: out <= 12'hf76;
      20'h065a5: out <= 12'hf76;
      20'h065a6: out <= 12'hf76;
      20'h065a7: out <= 12'hf76;
      20'h065a8: out <= 12'hfa9;
      20'h065a9: out <= 12'hfa9;
      20'h065aa: out <= 12'hfa9;
      20'h065ab: out <= 12'hfa9;
      20'h065ac: out <= 12'hfa9;
      20'h065ad: out <= 12'hfa9;
      20'h065ae: out <= 12'hfa9;
      20'h065af: out <= 12'hfa9;
      20'h065b0: out <= 12'h000;
      20'h065b1: out <= 12'h000;
      20'h065b2: out <= 12'h000;
      20'h065b3: out <= 12'h000;
      20'h065b4: out <= 12'h000;
      20'h065b5: out <= 12'h000;
      20'h065b6: out <= 12'h000;
      20'h065b7: out <= 12'h000;
      20'h065b8: out <= 12'h000;
      20'h065b9: out <= 12'h000;
      20'h065ba: out <= 12'h000;
      20'h065bb: out <= 12'h000;
      20'h065bc: out <= 12'h000;
      20'h065bd: out <= 12'h000;
      20'h065be: out <= 12'h000;
      20'h065bf: out <= 12'h000;
      20'h065c0: out <= 12'h000;
      20'h065c1: out <= 12'h000;
      20'h065c2: out <= 12'h000;
      20'h065c3: out <= 12'h000;
      20'h065c4: out <= 12'h000;
      20'h065c5: out <= 12'h000;
      20'h065c6: out <= 12'h000;
      20'h065c7: out <= 12'h000;
      20'h065c8: out <= 12'h222;
      20'h065c9: out <= 12'h222;
      20'h065ca: out <= 12'h222;
      20'h065cb: out <= 12'h222;
      20'h065cc: out <= 12'h222;
      20'h065cd: out <= 12'h222;
      20'h065ce: out <= 12'h222;
      20'h065cf: out <= 12'h222;
      20'h065d0: out <= 12'h222;
      20'h065d1: out <= 12'h222;
      20'h065d2: out <= 12'h222;
      20'h065d3: out <= 12'h222;
      20'h065d4: out <= 12'h222;
      20'h065d5: out <= 12'h222;
      20'h065d6: out <= 12'h222;
      20'h065d7: out <= 12'h222;
      20'h065d8: out <= 12'h000;
      20'h065d9: out <= 12'h000;
      20'h065da: out <= 12'h000;
      20'h065db: out <= 12'h000;
      20'h065dc: out <= 12'h000;
      20'h065dd: out <= 12'h666;
      20'h065de: out <= 12'hbbb;
      20'h065df: out <= 12'hbbb;
      20'h065e0: out <= 12'hbbb;
      20'h065e1: out <= 12'hbbb;
      20'h065e2: out <= 12'hbbb;
      20'h065e3: out <= 12'h666;
      20'h065e4: out <= 12'h000;
      20'h065e5: out <= 12'h000;
      20'h065e6: out <= 12'h000;
      20'h065e7: out <= 12'h000;
      20'h065e8: out <= 12'h222;
      20'h065e9: out <= 12'h222;
      20'h065ea: out <= 12'h222;
      20'h065eb: out <= 12'h222;
      20'h065ec: out <= 12'h222;
      20'h065ed: out <= 12'h666;
      20'h065ee: out <= 12'hbbb;
      20'h065ef: out <= 12'hbbb;
      20'h065f0: out <= 12'hbbb;
      20'h065f1: out <= 12'hbbb;
      20'h065f2: out <= 12'hbbb;
      20'h065f3: out <= 12'h666;
      20'h065f4: out <= 12'h222;
      20'h065f5: out <= 12'h222;
      20'h065f6: out <= 12'h222;
      20'h065f7: out <= 12'h222;
      20'h065f8: out <= 12'h000;
      20'h065f9: out <= 12'h000;
      20'h065fa: out <= 12'h000;
      20'h065fb: out <= 12'h000;
      20'h065fc: out <= 12'h000;
      20'h065fd: out <= 12'h000;
      20'h065fe: out <= 12'h000;
      20'h065ff: out <= 12'h000;
      20'h06600: out <= 12'h000;
      20'h06601: out <= 12'h000;
      20'h06602: out <= 12'h000;
      20'h06603: out <= 12'h000;
      20'h06604: out <= 12'h000;
      20'h06605: out <= 12'h000;
      20'h06606: out <= 12'h000;
      20'h06607: out <= 12'h000;
      20'h06608: out <= 12'h222;
      20'h06609: out <= 12'h222;
      20'h0660a: out <= 12'h222;
      20'h0660b: out <= 12'h222;
      20'h0660c: out <= 12'h222;
      20'h0660d: out <= 12'h222;
      20'h0660e: out <= 12'h222;
      20'h0660f: out <= 12'h222;
      20'h06610: out <= 12'h222;
      20'h06611: out <= 12'h222;
      20'h06612: out <= 12'h222;
      20'h06613: out <= 12'h222;
      20'h06614: out <= 12'h222;
      20'h06615: out <= 12'h222;
      20'h06616: out <= 12'h222;
      20'h06617: out <= 12'h222;
      20'h06618: out <= 12'h000;
      20'h06619: out <= 12'h000;
      20'h0661a: out <= 12'h000;
      20'h0661b: out <= 12'h000;
      20'h0661c: out <= 12'h000;
      20'h0661d: out <= 12'h000;
      20'h0661e: out <= 12'h000;
      20'h0661f: out <= 12'h666;
      20'h06620: out <= 12'hfff;
      20'h06621: out <= 12'h666;
      20'h06622: out <= 12'h000;
      20'h06623: out <= 12'h000;
      20'h06624: out <= 12'h000;
      20'h06625: out <= 12'h000;
      20'h06626: out <= 12'h000;
      20'h06627: out <= 12'h000;
      20'h06628: out <= 12'h222;
      20'h06629: out <= 12'h222;
      20'h0662a: out <= 12'h222;
      20'h0662b: out <= 12'h222;
      20'h0662c: out <= 12'h222;
      20'h0662d: out <= 12'h222;
      20'h0662e: out <= 12'h222;
      20'h0662f: out <= 12'h666;
      20'h06630: out <= 12'hfff;
      20'h06631: out <= 12'h666;
      20'h06632: out <= 12'h222;
      20'h06633: out <= 12'h222;
      20'h06634: out <= 12'h222;
      20'h06635: out <= 12'h222;
      20'h06636: out <= 12'h222;
      20'h06637: out <= 12'h222;
      20'h06638: out <= 12'h603;
      20'h06639: out <= 12'h603;
      20'h0663a: out <= 12'h603;
      20'h0663b: out <= 12'h603;
      20'h0663c: out <= 12'h603;
      20'h0663d: out <= 12'h603;
      20'h0663e: out <= 12'h603;
      20'h0663f: out <= 12'h603;
      20'h06640: out <= 12'h603;
      20'h06641: out <= 12'h603;
      20'h06642: out <= 12'h603;
      20'h06643: out <= 12'h603;
      20'h06644: out <= 12'h603;
      20'h06645: out <= 12'h603;
      20'h06646: out <= 12'h603;
      20'h06647: out <= 12'h603;
      20'h06648: out <= 12'h603;
      20'h06649: out <= 12'h603;
      20'h0664a: out <= 12'h603;
      20'h0664b: out <= 12'h603;
      20'h0664c: out <= 12'h603;
      20'h0664d: out <= 12'h603;
      20'h0664e: out <= 12'h603;
      20'h0664f: out <= 12'h603;
      20'h06650: out <= 12'h603;
      20'h06651: out <= 12'h603;
      20'h06652: out <= 12'h603;
      20'h06653: out <= 12'h603;
      20'h06654: out <= 12'h603;
      20'h06655: out <= 12'h603;
      20'h06656: out <= 12'h603;
      20'h06657: out <= 12'h603;
      20'h06658: out <= 12'h603;
      20'h06659: out <= 12'h603;
      20'h0665a: out <= 12'h603;
      20'h0665b: out <= 12'h603;
      20'h0665c: out <= 12'h603;
      20'h0665d: out <= 12'h603;
      20'h0665e: out <= 12'h603;
      20'h0665f: out <= 12'h603;
      20'h06660: out <= 12'h603;
      20'h06661: out <= 12'h603;
      20'h06662: out <= 12'h603;
      20'h06663: out <= 12'h603;
      20'h06664: out <= 12'h603;
      20'h06665: out <= 12'h603;
      20'h06666: out <= 12'h603;
      20'h06667: out <= 12'h603;
      20'h06668: out <= 12'h603;
      20'h06669: out <= 12'h603;
      20'h0666a: out <= 12'h603;
      20'h0666b: out <= 12'h603;
      20'h0666c: out <= 12'h603;
      20'h0666d: out <= 12'h603;
      20'h0666e: out <= 12'h603;
      20'h0666f: out <= 12'h603;
      20'h06670: out <= 12'h603;
      20'h06671: out <= 12'h603;
      20'h06672: out <= 12'h603;
      20'h06673: out <= 12'h603;
      20'h06674: out <= 12'h603;
      20'h06675: out <= 12'h603;
      20'h06676: out <= 12'h603;
      20'h06677: out <= 12'h603;
      20'h06678: out <= 12'h603;
      20'h06679: out <= 12'h603;
      20'h0667a: out <= 12'h603;
      20'h0667b: out <= 12'h603;
      20'h0667c: out <= 12'h603;
      20'h0667d: out <= 12'h603;
      20'h0667e: out <= 12'h603;
      20'h0667f: out <= 12'h603;
      20'h06680: out <= 12'h603;
      20'h06681: out <= 12'h603;
      20'h06682: out <= 12'h603;
      20'h06683: out <= 12'h603;
      20'h06684: out <= 12'h603;
      20'h06685: out <= 12'h603;
      20'h06686: out <= 12'h603;
      20'h06687: out <= 12'h603;
      20'h06688: out <= 12'h603;
      20'h06689: out <= 12'h603;
      20'h0668a: out <= 12'h603;
      20'h0668b: out <= 12'h603;
      20'h0668c: out <= 12'h603;
      20'h0668d: out <= 12'h603;
      20'h0668e: out <= 12'h603;
      20'h0668f: out <= 12'h603;
      20'h06690: out <= 12'hee9;
      20'h06691: out <= 12'hf87;
      20'h06692: out <= 12'hee9;
      20'h06693: out <= 12'hb27;
      20'h06694: out <= 12'hb27;
      20'h06695: out <= 12'hb27;
      20'h06696: out <= 12'hf87;
      20'h06697: out <= 12'hb27;
      20'h06698: out <= 12'h000;
      20'h06699: out <= 12'h000;
      20'h0669a: out <= 12'h000;
      20'h0669b: out <= 12'h000;
      20'h0669c: out <= 12'h000;
      20'h0669d: out <= 12'h000;
      20'h0669e: out <= 12'h000;
      20'h0669f: out <= 12'h000;
      20'h066a0: out <= 12'hfa9;
      20'h066a1: out <= 12'hfa9;
      20'h066a2: out <= 12'hfa9;
      20'h066a3: out <= 12'hfa9;
      20'h066a4: out <= 12'hfa9;
      20'h066a5: out <= 12'hfa9;
      20'h066a6: out <= 12'hfa9;
      20'h066a7: out <= 12'hfa9;
      20'h066a8: out <= 12'hf76;
      20'h066a9: out <= 12'hf76;
      20'h066aa: out <= 12'hf76;
      20'h066ab: out <= 12'hf76;
      20'h066ac: out <= 12'hf76;
      20'h066ad: out <= 12'hf76;
      20'h066ae: out <= 12'hf76;
      20'h066af: out <= 12'hf76;
      20'h066b0: out <= 12'hfa9;
      20'h066b1: out <= 12'hfa9;
      20'h066b2: out <= 12'hfa9;
      20'h066b3: out <= 12'hfa9;
      20'h066b4: out <= 12'hfa9;
      20'h066b5: out <= 12'hfa9;
      20'h066b6: out <= 12'hfa9;
      20'h066b7: out <= 12'hfa9;
      20'h066b8: out <= 12'hf76;
      20'h066b9: out <= 12'hf76;
      20'h066ba: out <= 12'hf76;
      20'h066bb: out <= 12'hf76;
      20'h066bc: out <= 12'hf76;
      20'h066bd: out <= 12'hf76;
      20'h066be: out <= 12'hf76;
      20'h066bf: out <= 12'hf76;
      20'h066c0: out <= 12'hfa9;
      20'h066c1: out <= 12'hfa9;
      20'h066c2: out <= 12'hfa9;
      20'h066c3: out <= 12'hfa9;
      20'h066c4: out <= 12'hfa9;
      20'h066c5: out <= 12'hfa9;
      20'h066c6: out <= 12'hfa9;
      20'h066c7: out <= 12'hfa9;
      20'h066c8: out <= 12'h000;
      20'h066c9: out <= 12'h000;
      20'h066ca: out <= 12'h000;
      20'h066cb: out <= 12'h000;
      20'h066cc: out <= 12'h000;
      20'h066cd: out <= 12'h000;
      20'h066ce: out <= 12'h000;
      20'h066cf: out <= 12'h000;
      20'h066d0: out <= 12'h000;
      20'h066d1: out <= 12'h000;
      20'h066d2: out <= 12'h000;
      20'h066d3: out <= 12'h000;
      20'h066d4: out <= 12'h000;
      20'h066d5: out <= 12'h000;
      20'h066d6: out <= 12'h000;
      20'h066d7: out <= 12'h000;
      20'h066d8: out <= 12'h000;
      20'h066d9: out <= 12'h000;
      20'h066da: out <= 12'h000;
      20'h066db: out <= 12'h000;
      20'h066dc: out <= 12'h000;
      20'h066dd: out <= 12'h000;
      20'h066de: out <= 12'h000;
      20'h066df: out <= 12'h000;
      20'h066e0: out <= 12'h222;
      20'h066e1: out <= 12'h222;
      20'h066e2: out <= 12'h222;
      20'h066e3: out <= 12'h222;
      20'h066e4: out <= 12'h222;
      20'h066e5: out <= 12'h222;
      20'h066e6: out <= 12'h222;
      20'h066e7: out <= 12'h222;
      20'h066e8: out <= 12'h222;
      20'h066e9: out <= 12'h222;
      20'h066ea: out <= 12'h222;
      20'h066eb: out <= 12'h222;
      20'h066ec: out <= 12'h222;
      20'h066ed: out <= 12'h222;
      20'h066ee: out <= 12'h222;
      20'h066ef: out <= 12'h222;
      20'h066f0: out <= 12'h000;
      20'h066f1: out <= 12'h000;
      20'h066f2: out <= 12'h000;
      20'h066f3: out <= 12'h000;
      20'h066f4: out <= 12'h000;
      20'h066f5: out <= 12'h000;
      20'h066f6: out <= 12'h666;
      20'h066f7: out <= 12'h666;
      20'h066f8: out <= 12'h666;
      20'h066f9: out <= 12'h666;
      20'h066fa: out <= 12'h666;
      20'h066fb: out <= 12'h000;
      20'h066fc: out <= 12'h000;
      20'h066fd: out <= 12'h000;
      20'h066fe: out <= 12'h000;
      20'h066ff: out <= 12'h000;
      20'h06700: out <= 12'h222;
      20'h06701: out <= 12'h222;
      20'h06702: out <= 12'h222;
      20'h06703: out <= 12'h222;
      20'h06704: out <= 12'h222;
      20'h06705: out <= 12'h222;
      20'h06706: out <= 12'h666;
      20'h06707: out <= 12'h666;
      20'h06708: out <= 12'h666;
      20'h06709: out <= 12'h666;
      20'h0670a: out <= 12'h666;
      20'h0670b: out <= 12'h222;
      20'h0670c: out <= 12'h222;
      20'h0670d: out <= 12'h222;
      20'h0670e: out <= 12'h222;
      20'h0670f: out <= 12'h222;
      20'h06710: out <= 12'h000;
      20'h06711: out <= 12'h000;
      20'h06712: out <= 12'h000;
      20'h06713: out <= 12'h000;
      20'h06714: out <= 12'h000;
      20'h06715: out <= 12'h000;
      20'h06716: out <= 12'h000;
      20'h06717: out <= 12'h000;
      20'h06718: out <= 12'h000;
      20'h06719: out <= 12'h000;
      20'h0671a: out <= 12'h000;
      20'h0671b: out <= 12'h000;
      20'h0671c: out <= 12'h000;
      20'h0671d: out <= 12'h000;
      20'h0671e: out <= 12'h000;
      20'h0671f: out <= 12'h000;
      20'h06720: out <= 12'h222;
      20'h06721: out <= 12'h222;
      20'h06722: out <= 12'h222;
      20'h06723: out <= 12'h222;
      20'h06724: out <= 12'h222;
      20'h06725: out <= 12'h222;
      20'h06726: out <= 12'h222;
      20'h06727: out <= 12'h222;
      20'h06728: out <= 12'h222;
      20'h06729: out <= 12'h222;
      20'h0672a: out <= 12'h222;
      20'h0672b: out <= 12'h222;
      20'h0672c: out <= 12'h222;
      20'h0672d: out <= 12'h222;
      20'h0672e: out <= 12'h222;
      20'h0672f: out <= 12'h222;
      20'h06730: out <= 12'h000;
      20'h06731: out <= 12'h000;
      20'h06732: out <= 12'h000;
      20'h06733: out <= 12'h000;
      20'h06734: out <= 12'h000;
      20'h06735: out <= 12'h000;
      20'h06736: out <= 12'h000;
      20'h06737: out <= 12'h666;
      20'h06738: out <= 12'hfff;
      20'h06739: out <= 12'h666;
      20'h0673a: out <= 12'h000;
      20'h0673b: out <= 12'h000;
      20'h0673c: out <= 12'h000;
      20'h0673d: out <= 12'h000;
      20'h0673e: out <= 12'h000;
      20'h0673f: out <= 12'h000;
      20'h06740: out <= 12'h222;
      20'h06741: out <= 12'h222;
      20'h06742: out <= 12'h222;
      20'h06743: out <= 12'h222;
      20'h06744: out <= 12'h222;
      20'h06745: out <= 12'h222;
      20'h06746: out <= 12'h222;
      20'h06747: out <= 12'h666;
      20'h06748: out <= 12'hfff;
      20'h06749: out <= 12'h666;
      20'h0674a: out <= 12'h222;
      20'h0674b: out <= 12'h222;
      20'h0674c: out <= 12'h222;
      20'h0674d: out <= 12'h222;
      20'h0674e: out <= 12'h222;
      20'h0674f: out <= 12'h222;
      20'h06750: out <= 12'h603;
      20'h06751: out <= 12'h603;
      20'h06752: out <= 12'h603;
      20'h06753: out <= 12'h603;
      20'h06754: out <= 12'h603;
      20'h06755: out <= 12'h603;
      20'h06756: out <= 12'h603;
      20'h06757: out <= 12'h603;
      20'h06758: out <= 12'h603;
      20'h06759: out <= 12'h603;
      20'h0675a: out <= 12'h603;
      20'h0675b: out <= 12'h603;
      20'h0675c: out <= 12'h603;
      20'h0675d: out <= 12'h603;
      20'h0675e: out <= 12'h603;
      20'h0675f: out <= 12'h603;
      20'h06760: out <= 12'h603;
      20'h06761: out <= 12'h603;
      20'h06762: out <= 12'h603;
      20'h06763: out <= 12'h603;
      20'h06764: out <= 12'h603;
      20'h06765: out <= 12'h603;
      20'h06766: out <= 12'h603;
      20'h06767: out <= 12'h603;
      20'h06768: out <= 12'h603;
      20'h06769: out <= 12'h603;
      20'h0676a: out <= 12'h603;
      20'h0676b: out <= 12'h603;
      20'h0676c: out <= 12'h603;
      20'h0676d: out <= 12'h603;
      20'h0676e: out <= 12'h603;
      20'h0676f: out <= 12'h603;
      20'h06770: out <= 12'h603;
      20'h06771: out <= 12'h603;
      20'h06772: out <= 12'h603;
      20'h06773: out <= 12'h603;
      20'h06774: out <= 12'h603;
      20'h06775: out <= 12'h603;
      20'h06776: out <= 12'h603;
      20'h06777: out <= 12'h603;
      20'h06778: out <= 12'h603;
      20'h06779: out <= 12'h603;
      20'h0677a: out <= 12'h603;
      20'h0677b: out <= 12'h603;
      20'h0677c: out <= 12'h603;
      20'h0677d: out <= 12'h603;
      20'h0677e: out <= 12'h603;
      20'h0677f: out <= 12'h603;
      20'h06780: out <= 12'h603;
      20'h06781: out <= 12'h603;
      20'h06782: out <= 12'h603;
      20'h06783: out <= 12'h603;
      20'h06784: out <= 12'h603;
      20'h06785: out <= 12'h603;
      20'h06786: out <= 12'h603;
      20'h06787: out <= 12'h603;
      20'h06788: out <= 12'h603;
      20'h06789: out <= 12'h603;
      20'h0678a: out <= 12'h603;
      20'h0678b: out <= 12'h603;
      20'h0678c: out <= 12'h603;
      20'h0678d: out <= 12'h603;
      20'h0678e: out <= 12'h603;
      20'h0678f: out <= 12'h603;
      20'h06790: out <= 12'h603;
      20'h06791: out <= 12'h603;
      20'h06792: out <= 12'h603;
      20'h06793: out <= 12'h603;
      20'h06794: out <= 12'h603;
      20'h06795: out <= 12'h603;
      20'h06796: out <= 12'h603;
      20'h06797: out <= 12'h603;
      20'h06798: out <= 12'h603;
      20'h06799: out <= 12'h603;
      20'h0679a: out <= 12'h603;
      20'h0679b: out <= 12'h603;
      20'h0679c: out <= 12'h603;
      20'h0679d: out <= 12'h603;
      20'h0679e: out <= 12'h603;
      20'h0679f: out <= 12'h603;
      20'h067a0: out <= 12'h603;
      20'h067a1: out <= 12'h603;
      20'h067a2: out <= 12'h603;
      20'h067a3: out <= 12'h603;
      20'h067a4: out <= 12'h603;
      20'h067a5: out <= 12'h603;
      20'h067a6: out <= 12'h603;
      20'h067a7: out <= 12'h603;
      20'h067a8: out <= 12'hee9;
      20'h067a9: out <= 12'hf87;
      20'h067aa: out <= 12'hf87;
      20'h067ab: out <= 12'hf87;
      20'h067ac: out <= 12'hf87;
      20'h067ad: out <= 12'hf87;
      20'h067ae: out <= 12'hf87;
      20'h067af: out <= 12'hb27;
      20'h067b0: out <= 12'h000;
      20'h067b1: out <= 12'h000;
      20'h067b2: out <= 12'h000;
      20'h067b3: out <= 12'h000;
      20'h067b4: out <= 12'h000;
      20'h067b5: out <= 12'h000;
      20'h067b6: out <= 12'h000;
      20'h067b7: out <= 12'h000;
      20'h067b8: out <= 12'hfa9;
      20'h067b9: out <= 12'hfa9;
      20'h067ba: out <= 12'hfa9;
      20'h067bb: out <= 12'hfa9;
      20'h067bc: out <= 12'hfa9;
      20'h067bd: out <= 12'hfa9;
      20'h067be: out <= 12'hfa9;
      20'h067bf: out <= 12'hfa9;
      20'h067c0: out <= 12'hf76;
      20'h067c1: out <= 12'hf76;
      20'h067c2: out <= 12'hf76;
      20'h067c3: out <= 12'hf76;
      20'h067c4: out <= 12'hf76;
      20'h067c5: out <= 12'hf76;
      20'h067c6: out <= 12'hf76;
      20'h067c7: out <= 12'hf76;
      20'h067c8: out <= 12'hfa9;
      20'h067c9: out <= 12'hfa9;
      20'h067ca: out <= 12'hfa9;
      20'h067cb: out <= 12'hfa9;
      20'h067cc: out <= 12'hfa9;
      20'h067cd: out <= 12'hfa9;
      20'h067ce: out <= 12'hfa9;
      20'h067cf: out <= 12'hfa9;
      20'h067d0: out <= 12'hf76;
      20'h067d1: out <= 12'hf76;
      20'h067d2: out <= 12'hf76;
      20'h067d3: out <= 12'hf76;
      20'h067d4: out <= 12'hf76;
      20'h067d5: out <= 12'hf76;
      20'h067d6: out <= 12'hf76;
      20'h067d7: out <= 12'hf76;
      20'h067d8: out <= 12'hfa9;
      20'h067d9: out <= 12'hfa9;
      20'h067da: out <= 12'hfa9;
      20'h067db: out <= 12'hfa9;
      20'h067dc: out <= 12'hfa9;
      20'h067dd: out <= 12'hfa9;
      20'h067de: out <= 12'hfa9;
      20'h067df: out <= 12'hfa9;
      20'h067e0: out <= 12'h000;
      20'h067e1: out <= 12'h000;
      20'h067e2: out <= 12'h000;
      20'h067e3: out <= 12'h000;
      20'h067e4: out <= 12'h000;
      20'h067e5: out <= 12'h000;
      20'h067e6: out <= 12'h000;
      20'h067e7: out <= 12'h000;
      20'h067e8: out <= 12'h000;
      20'h067e9: out <= 12'h000;
      20'h067ea: out <= 12'h000;
      20'h067eb: out <= 12'h000;
      20'h067ec: out <= 12'h000;
      20'h067ed: out <= 12'h000;
      20'h067ee: out <= 12'h000;
      20'h067ef: out <= 12'h000;
      20'h067f0: out <= 12'h000;
      20'h067f1: out <= 12'h000;
      20'h067f2: out <= 12'h000;
      20'h067f3: out <= 12'h000;
      20'h067f4: out <= 12'h000;
      20'h067f5: out <= 12'h000;
      20'h067f6: out <= 12'h000;
      20'h067f7: out <= 12'h000;
      20'h067f8: out <= 12'h222;
      20'h067f9: out <= 12'h222;
      20'h067fa: out <= 12'h222;
      20'h067fb: out <= 12'h222;
      20'h067fc: out <= 12'h222;
      20'h067fd: out <= 12'h222;
      20'h067fe: out <= 12'h222;
      20'h067ff: out <= 12'h222;
      20'h06800: out <= 12'h222;
      20'h06801: out <= 12'h222;
      20'h06802: out <= 12'h222;
      20'h06803: out <= 12'h222;
      20'h06804: out <= 12'h222;
      20'h06805: out <= 12'h222;
      20'h06806: out <= 12'h222;
      20'h06807: out <= 12'h222;
      20'h06808: out <= 12'h000;
      20'h06809: out <= 12'h000;
      20'h0680a: out <= 12'h000;
      20'h0680b: out <= 12'h000;
      20'h0680c: out <= 12'h000;
      20'h0680d: out <= 12'h000;
      20'h0680e: out <= 12'h000;
      20'h0680f: out <= 12'h000;
      20'h06810: out <= 12'h000;
      20'h06811: out <= 12'h000;
      20'h06812: out <= 12'h000;
      20'h06813: out <= 12'h000;
      20'h06814: out <= 12'h000;
      20'h06815: out <= 12'h000;
      20'h06816: out <= 12'h000;
      20'h06817: out <= 12'h000;
      20'h06818: out <= 12'h222;
      20'h06819: out <= 12'h222;
      20'h0681a: out <= 12'h222;
      20'h0681b: out <= 12'h222;
      20'h0681c: out <= 12'h222;
      20'h0681d: out <= 12'h222;
      20'h0681e: out <= 12'h222;
      20'h0681f: out <= 12'h222;
      20'h06820: out <= 12'h222;
      20'h06821: out <= 12'h222;
      20'h06822: out <= 12'h222;
      20'h06823: out <= 12'h222;
      20'h06824: out <= 12'h222;
      20'h06825: out <= 12'h222;
      20'h06826: out <= 12'h222;
      20'h06827: out <= 12'h222;
      20'h06828: out <= 12'h000;
      20'h06829: out <= 12'h000;
      20'h0682a: out <= 12'h000;
      20'h0682b: out <= 12'h000;
      20'h0682c: out <= 12'h000;
      20'h0682d: out <= 12'h000;
      20'h0682e: out <= 12'h000;
      20'h0682f: out <= 12'h000;
      20'h06830: out <= 12'h000;
      20'h06831: out <= 12'h000;
      20'h06832: out <= 12'h000;
      20'h06833: out <= 12'h000;
      20'h06834: out <= 12'h000;
      20'h06835: out <= 12'h000;
      20'h06836: out <= 12'h000;
      20'h06837: out <= 12'h000;
      20'h06838: out <= 12'h222;
      20'h06839: out <= 12'h222;
      20'h0683a: out <= 12'h222;
      20'h0683b: out <= 12'h222;
      20'h0683c: out <= 12'h222;
      20'h0683d: out <= 12'h222;
      20'h0683e: out <= 12'h222;
      20'h0683f: out <= 12'h222;
      20'h06840: out <= 12'h222;
      20'h06841: out <= 12'h222;
      20'h06842: out <= 12'h222;
      20'h06843: out <= 12'h222;
      20'h06844: out <= 12'h222;
      20'h06845: out <= 12'h222;
      20'h06846: out <= 12'h222;
      20'h06847: out <= 12'h222;
      20'h06848: out <= 12'h000;
      20'h06849: out <= 12'h000;
      20'h0684a: out <= 12'h000;
      20'h0684b: out <= 12'h000;
      20'h0684c: out <= 12'h000;
      20'h0684d: out <= 12'h000;
      20'h0684e: out <= 12'h000;
      20'h0684f: out <= 12'h666;
      20'h06850: out <= 12'hfff;
      20'h06851: out <= 12'h666;
      20'h06852: out <= 12'h000;
      20'h06853: out <= 12'h000;
      20'h06854: out <= 12'h000;
      20'h06855: out <= 12'h000;
      20'h06856: out <= 12'h000;
      20'h06857: out <= 12'h000;
      20'h06858: out <= 12'h222;
      20'h06859: out <= 12'h222;
      20'h0685a: out <= 12'h222;
      20'h0685b: out <= 12'h222;
      20'h0685c: out <= 12'h222;
      20'h0685d: out <= 12'h222;
      20'h0685e: out <= 12'h222;
      20'h0685f: out <= 12'h666;
      20'h06860: out <= 12'hfff;
      20'h06861: out <= 12'h666;
      20'h06862: out <= 12'h222;
      20'h06863: out <= 12'h222;
      20'h06864: out <= 12'h222;
      20'h06865: out <= 12'h222;
      20'h06866: out <= 12'h222;
      20'h06867: out <= 12'h222;
      20'h06868: out <= 12'h603;
      20'h06869: out <= 12'h603;
      20'h0686a: out <= 12'h603;
      20'h0686b: out <= 12'h603;
      20'h0686c: out <= 12'h603;
      20'h0686d: out <= 12'h603;
      20'h0686e: out <= 12'h603;
      20'h0686f: out <= 12'h603;
      20'h06870: out <= 12'h603;
      20'h06871: out <= 12'h603;
      20'h06872: out <= 12'h603;
      20'h06873: out <= 12'h603;
      20'h06874: out <= 12'h603;
      20'h06875: out <= 12'h603;
      20'h06876: out <= 12'h603;
      20'h06877: out <= 12'h603;
      20'h06878: out <= 12'h603;
      20'h06879: out <= 12'h603;
      20'h0687a: out <= 12'h603;
      20'h0687b: out <= 12'h603;
      20'h0687c: out <= 12'h603;
      20'h0687d: out <= 12'h603;
      20'h0687e: out <= 12'h603;
      20'h0687f: out <= 12'h603;
      20'h06880: out <= 12'h603;
      20'h06881: out <= 12'h603;
      20'h06882: out <= 12'h603;
      20'h06883: out <= 12'h603;
      20'h06884: out <= 12'h603;
      20'h06885: out <= 12'h603;
      20'h06886: out <= 12'h603;
      20'h06887: out <= 12'h603;
      20'h06888: out <= 12'h603;
      20'h06889: out <= 12'h603;
      20'h0688a: out <= 12'h603;
      20'h0688b: out <= 12'h603;
      20'h0688c: out <= 12'h603;
      20'h0688d: out <= 12'h603;
      20'h0688e: out <= 12'h603;
      20'h0688f: out <= 12'h603;
      20'h06890: out <= 12'h603;
      20'h06891: out <= 12'h603;
      20'h06892: out <= 12'h603;
      20'h06893: out <= 12'h603;
      20'h06894: out <= 12'h603;
      20'h06895: out <= 12'h603;
      20'h06896: out <= 12'h603;
      20'h06897: out <= 12'h603;
      20'h06898: out <= 12'h603;
      20'h06899: out <= 12'h603;
      20'h0689a: out <= 12'h603;
      20'h0689b: out <= 12'h603;
      20'h0689c: out <= 12'h603;
      20'h0689d: out <= 12'h603;
      20'h0689e: out <= 12'h603;
      20'h0689f: out <= 12'h603;
      20'h068a0: out <= 12'h603;
      20'h068a1: out <= 12'h603;
      20'h068a2: out <= 12'h603;
      20'h068a3: out <= 12'h603;
      20'h068a4: out <= 12'h603;
      20'h068a5: out <= 12'h603;
      20'h068a6: out <= 12'h603;
      20'h068a7: out <= 12'h603;
      20'h068a8: out <= 12'h603;
      20'h068a9: out <= 12'h603;
      20'h068aa: out <= 12'h603;
      20'h068ab: out <= 12'h603;
      20'h068ac: out <= 12'h603;
      20'h068ad: out <= 12'h603;
      20'h068ae: out <= 12'h603;
      20'h068af: out <= 12'h603;
      20'h068b0: out <= 12'h603;
      20'h068b1: out <= 12'h603;
      20'h068b2: out <= 12'h603;
      20'h068b3: out <= 12'h603;
      20'h068b4: out <= 12'h603;
      20'h068b5: out <= 12'h603;
      20'h068b6: out <= 12'h603;
      20'h068b7: out <= 12'h603;
      20'h068b8: out <= 12'h603;
      20'h068b9: out <= 12'h603;
      20'h068ba: out <= 12'h603;
      20'h068bb: out <= 12'h603;
      20'h068bc: out <= 12'h603;
      20'h068bd: out <= 12'h603;
      20'h068be: out <= 12'h603;
      20'h068bf: out <= 12'h603;
      20'h068c0: out <= 12'hb27;
      20'h068c1: out <= 12'hb27;
      20'h068c2: out <= 12'hb27;
      20'h068c3: out <= 12'hb27;
      20'h068c4: out <= 12'hb27;
      20'h068c5: out <= 12'hb27;
      20'h068c6: out <= 12'hb27;
      20'h068c7: out <= 12'hb27;
      20'h068c8: out <= 12'h000;
      20'h068c9: out <= 12'h000;
      20'h068ca: out <= 12'h000;
      20'h068cb: out <= 12'h000;
      20'h068cc: out <= 12'h000;
      20'h068cd: out <= 12'h000;
      20'h068ce: out <= 12'h000;
      20'h068cf: out <= 12'h000;
      20'h068d0: out <= 12'hfa9;
      20'h068d1: out <= 12'hfa9;
      20'h068d2: out <= 12'hfa9;
      20'h068d3: out <= 12'hfa9;
      20'h068d4: out <= 12'hfa9;
      20'h068d5: out <= 12'hfa9;
      20'h068d6: out <= 12'hfa9;
      20'h068d7: out <= 12'hfa9;
      20'h068d8: out <= 12'hf76;
      20'h068d9: out <= 12'hf76;
      20'h068da: out <= 12'hf76;
      20'h068db: out <= 12'hf76;
      20'h068dc: out <= 12'hf76;
      20'h068dd: out <= 12'hf76;
      20'h068de: out <= 12'hf76;
      20'h068df: out <= 12'hf76;
      20'h068e0: out <= 12'hfa9;
      20'h068e1: out <= 12'hfa9;
      20'h068e2: out <= 12'hfa9;
      20'h068e3: out <= 12'hfa9;
      20'h068e4: out <= 12'hfa9;
      20'h068e5: out <= 12'hfa9;
      20'h068e6: out <= 12'hfa9;
      20'h068e7: out <= 12'hfa9;
      20'h068e8: out <= 12'hf76;
      20'h068e9: out <= 12'hf76;
      20'h068ea: out <= 12'hf76;
      20'h068eb: out <= 12'hf76;
      20'h068ec: out <= 12'hf76;
      20'h068ed: out <= 12'hf76;
      20'h068ee: out <= 12'hf76;
      20'h068ef: out <= 12'hf76;
      20'h068f0: out <= 12'hfa9;
      20'h068f1: out <= 12'hfa9;
      20'h068f2: out <= 12'hfa9;
      20'h068f3: out <= 12'hfa9;
      20'h068f4: out <= 12'hfa9;
      20'h068f5: out <= 12'hfa9;
      20'h068f6: out <= 12'hfa9;
      20'h068f7: out <= 12'hfa9;
      20'h068f8: out <= 12'h000;
      20'h068f9: out <= 12'h000;
      20'h068fa: out <= 12'h000;
      20'h068fb: out <= 12'h000;
      20'h068fc: out <= 12'h000;
      20'h068fd: out <= 12'h000;
      20'h068fe: out <= 12'h000;
      20'h068ff: out <= 12'h000;
      20'h06900: out <= 12'h222;
      20'h06901: out <= 12'h222;
      20'h06902: out <= 12'h222;
      20'h06903: out <= 12'h222;
      20'h06904: out <= 12'h222;
      20'h06905: out <= 12'h222;
      20'h06906: out <= 12'h222;
      20'h06907: out <= 12'h222;
      20'h06908: out <= 12'h222;
      20'h06909: out <= 12'h222;
      20'h0690a: out <= 12'h222;
      20'h0690b: out <= 12'h222;
      20'h0690c: out <= 12'h222;
      20'h0690d: out <= 12'h222;
      20'h0690e: out <= 12'h222;
      20'h0690f: out <= 12'h222;
      20'h06910: out <= 12'h000;
      20'h06911: out <= 12'h000;
      20'h06912: out <= 12'h000;
      20'h06913: out <= 12'h000;
      20'h06914: out <= 12'h000;
      20'h06915: out <= 12'h000;
      20'h06916: out <= 12'h000;
      20'h06917: out <= 12'h000;
      20'h06918: out <= 12'h000;
      20'h06919: out <= 12'h000;
      20'h0691a: out <= 12'h000;
      20'h0691b: out <= 12'h000;
      20'h0691c: out <= 12'h000;
      20'h0691d: out <= 12'h000;
      20'h0691e: out <= 12'h000;
      20'h0691f: out <= 12'h000;
      20'h06920: out <= 12'h222;
      20'h06921: out <= 12'h222;
      20'h06922: out <= 12'h222;
      20'h06923: out <= 12'h222;
      20'h06924: out <= 12'h222;
      20'h06925: out <= 12'h222;
      20'h06926: out <= 12'h666;
      20'h06927: out <= 12'hbbb;
      20'h06928: out <= 12'hfff;
      20'h06929: out <= 12'hbbb;
      20'h0692a: out <= 12'h666;
      20'h0692b: out <= 12'h222;
      20'h0692c: out <= 12'h222;
      20'h0692d: out <= 12'h222;
      20'h0692e: out <= 12'h222;
      20'h0692f: out <= 12'h222;
      20'h06930: out <= 12'h000;
      20'h06931: out <= 12'h000;
      20'h06932: out <= 12'h000;
      20'h06933: out <= 12'h000;
      20'h06934: out <= 12'h000;
      20'h06935: out <= 12'h000;
      20'h06936: out <= 12'h666;
      20'h06937: out <= 12'hbbb;
      20'h06938: out <= 12'hfff;
      20'h06939: out <= 12'hbbb;
      20'h0693a: out <= 12'h666;
      20'h0693b: out <= 12'h000;
      20'h0693c: out <= 12'h000;
      20'h0693d: out <= 12'h000;
      20'h0693e: out <= 12'h000;
      20'h0693f: out <= 12'h000;
      20'h06940: out <= 12'h222;
      20'h06941: out <= 12'h222;
      20'h06942: out <= 12'h222;
      20'h06943: out <= 12'h222;
      20'h06944: out <= 12'h222;
      20'h06945: out <= 12'h222;
      20'h06946: out <= 12'h222;
      20'h06947: out <= 12'h222;
      20'h06948: out <= 12'h222;
      20'h06949: out <= 12'h222;
      20'h0694a: out <= 12'h222;
      20'h0694b: out <= 12'h222;
      20'h0694c: out <= 12'h222;
      20'h0694d: out <= 12'h222;
      20'h0694e: out <= 12'h222;
      20'h0694f: out <= 12'h222;
      20'h06950: out <= 12'h000;
      20'h06951: out <= 12'h000;
      20'h06952: out <= 12'h000;
      20'h06953: out <= 12'h000;
      20'h06954: out <= 12'h000;
      20'h06955: out <= 12'h000;
      20'h06956: out <= 12'h000;
      20'h06957: out <= 12'h000;
      20'h06958: out <= 12'h000;
      20'h06959: out <= 12'h000;
      20'h0695a: out <= 12'h000;
      20'h0695b: out <= 12'h000;
      20'h0695c: out <= 12'h000;
      20'h0695d: out <= 12'h000;
      20'h0695e: out <= 12'h000;
      20'h0695f: out <= 12'h000;
      20'h06960: out <= 12'h222;
      20'h06961: out <= 12'h222;
      20'h06962: out <= 12'h222;
      20'h06963: out <= 12'h222;
      20'h06964: out <= 12'h222;
      20'h06965: out <= 12'h222;
      20'h06966: out <= 12'h222;
      20'h06967: out <= 12'h222;
      20'h06968: out <= 12'h222;
      20'h06969: out <= 12'h222;
      20'h0696a: out <= 12'h222;
      20'h0696b: out <= 12'h222;
      20'h0696c: out <= 12'h222;
      20'h0696d: out <= 12'h222;
      20'h0696e: out <= 12'h222;
      20'h0696f: out <= 12'h222;
      20'h06970: out <= 12'h000;
      20'h06971: out <= 12'h000;
      20'h06972: out <= 12'h000;
      20'h06973: out <= 12'h000;
      20'h06974: out <= 12'h000;
      20'h06975: out <= 12'h000;
      20'h06976: out <= 12'h000;
      20'h06977: out <= 12'h000;
      20'h06978: out <= 12'h000;
      20'h06979: out <= 12'h000;
      20'h0697a: out <= 12'h000;
      20'h0697b: out <= 12'h000;
      20'h0697c: out <= 12'h000;
      20'h0697d: out <= 12'h000;
      20'h0697e: out <= 12'h000;
      20'h0697f: out <= 12'h000;
      20'h06980: out <= 12'h603;
      20'h06981: out <= 12'h603;
      20'h06982: out <= 12'h603;
      20'h06983: out <= 12'h603;
      20'h06984: out <= 12'h603;
      20'h06985: out <= 12'h603;
      20'h06986: out <= 12'h603;
      20'h06987: out <= 12'h603;
      20'h06988: out <= 12'h603;
      20'h06989: out <= 12'h603;
      20'h0698a: out <= 12'h603;
      20'h0698b: out <= 12'h603;
      20'h0698c: out <= 12'hee9;
      20'h0698d: out <= 12'hee9;
      20'h0698e: out <= 12'hee9;
      20'h0698f: out <= 12'hee9;
      20'h06990: out <= 12'hee9;
      20'h06991: out <= 12'hee9;
      20'h06992: out <= 12'hee9;
      20'h06993: out <= 12'hb27;
      20'h06994: out <= 12'hee9;
      20'h06995: out <= 12'hee9;
      20'h06996: out <= 12'hee9;
      20'h06997: out <= 12'hee9;
      20'h06998: out <= 12'hee9;
      20'h06999: out <= 12'hee9;
      20'h0699a: out <= 12'hee9;
      20'h0699b: out <= 12'hb27;
      20'h0699c: out <= 12'hee9;
      20'h0699d: out <= 12'hee9;
      20'h0699e: out <= 12'hee9;
      20'h0699f: out <= 12'hee9;
      20'h069a0: out <= 12'hee9;
      20'h069a1: out <= 12'hee9;
      20'h069a2: out <= 12'hee9;
      20'h069a3: out <= 12'hb27;
      20'h069a4: out <= 12'hee9;
      20'h069a5: out <= 12'hee9;
      20'h069a6: out <= 12'hee9;
      20'h069a7: out <= 12'hee9;
      20'h069a8: out <= 12'hee9;
      20'h069a9: out <= 12'hee9;
      20'h069aa: out <= 12'hee9;
      20'h069ab: out <= 12'hb27;
      20'h069ac: out <= 12'h603;
      20'h069ad: out <= 12'h603;
      20'h069ae: out <= 12'h603;
      20'h069af: out <= 12'h603;
      20'h069b0: out <= 12'h603;
      20'h069b1: out <= 12'h603;
      20'h069b2: out <= 12'h603;
      20'h069b3: out <= 12'h603;
      20'h069b4: out <= 12'h603;
      20'h069b5: out <= 12'h603;
      20'h069b6: out <= 12'h603;
      20'h069b7: out <= 12'h603;
      20'h069b8: out <= 12'h603;
      20'h069b9: out <= 12'h603;
      20'h069ba: out <= 12'h603;
      20'h069bb: out <= 12'h603;
      20'h069bc: out <= 12'h603;
      20'h069bd: out <= 12'h603;
      20'h069be: out <= 12'h603;
      20'h069bf: out <= 12'h603;
      20'h069c0: out <= 12'h603;
      20'h069c1: out <= 12'h603;
      20'h069c2: out <= 12'h603;
      20'h069c3: out <= 12'h603;
      20'h069c4: out <= 12'h603;
      20'h069c5: out <= 12'h603;
      20'h069c6: out <= 12'h603;
      20'h069c7: out <= 12'h603;
      20'h069c8: out <= 12'h603;
      20'h069c9: out <= 12'h603;
      20'h069ca: out <= 12'h603;
      20'h069cb: out <= 12'h603;
      20'h069cc: out <= 12'h603;
      20'h069cd: out <= 12'h603;
      20'h069ce: out <= 12'h603;
      20'h069cf: out <= 12'h603;
      20'h069d0: out <= 12'h603;
      20'h069d1: out <= 12'h603;
      20'h069d2: out <= 12'h603;
      20'h069d3: out <= 12'h603;
      20'h069d4: out <= 12'h603;
      20'h069d5: out <= 12'h603;
      20'h069d6: out <= 12'h603;
      20'h069d7: out <= 12'h603;
      20'h069d8: out <= 12'hee9;
      20'h069d9: out <= 12'hee9;
      20'h069da: out <= 12'hee9;
      20'h069db: out <= 12'hee9;
      20'h069dc: out <= 12'hee9;
      20'h069dd: out <= 12'hee9;
      20'h069de: out <= 12'hee9;
      20'h069df: out <= 12'hb27;
      20'h069e0: out <= 12'h000;
      20'h069e1: out <= 12'h000;
      20'h069e2: out <= 12'h000;
      20'h069e3: out <= 12'h000;
      20'h069e4: out <= 12'h000;
      20'h069e5: out <= 12'h000;
      20'h069e6: out <= 12'h000;
      20'h069e7: out <= 12'h000;
      20'h069e8: out <= 12'h777;
      20'h069e9: out <= 12'h777;
      20'h069ea: out <= 12'h777;
      20'h069eb: out <= 12'h777;
      20'h069ec: out <= 12'h777;
      20'h069ed: out <= 12'h777;
      20'h069ee: out <= 12'h777;
      20'h069ef: out <= 12'h777;
      20'h069f0: out <= 12'h777;
      20'h069f1: out <= 12'h777;
      20'h069f2: out <= 12'h777;
      20'h069f3: out <= 12'h777;
      20'h069f4: out <= 12'h777;
      20'h069f5: out <= 12'h777;
      20'h069f6: out <= 12'h777;
      20'h069f7: out <= 12'h777;
      20'h069f8: out <= 12'h000;
      20'h069f9: out <= 12'h000;
      20'h069fa: out <= 12'h000;
      20'h069fb: out <= 12'h000;
      20'h069fc: out <= 12'h000;
      20'h069fd: out <= 12'h000;
      20'h069fe: out <= 12'h000;
      20'h069ff: out <= 12'h000;
      20'h06a00: out <= 12'h000;
      20'h06a01: out <= 12'h000;
      20'h06a02: out <= 12'h000;
      20'h06a03: out <= 12'h000;
      20'h06a04: out <= 12'h000;
      20'h06a05: out <= 12'h000;
      20'h06a06: out <= 12'h000;
      20'h06a07: out <= 12'h000;
      20'h06a08: out <= 12'h000;
      20'h06a09: out <= 12'h000;
      20'h06a0a: out <= 12'h000;
      20'h06a0b: out <= 12'h000;
      20'h06a0c: out <= 12'h000;
      20'h06a0d: out <= 12'h000;
      20'h06a0e: out <= 12'h000;
      20'h06a0f: out <= 12'h000;
      20'h06a10: out <= 12'h000;
      20'h06a11: out <= 12'h000;
      20'h06a12: out <= 12'h000;
      20'h06a13: out <= 12'h000;
      20'h06a14: out <= 12'h000;
      20'h06a15: out <= 12'h000;
      20'h06a16: out <= 12'h000;
      20'h06a17: out <= 12'h000;
      20'h06a18: out <= 12'h222;
      20'h06a19: out <= 12'h222;
      20'h06a1a: out <= 12'h222;
      20'h06a1b: out <= 12'h666;
      20'h06a1c: out <= 12'h222;
      20'h06a1d: out <= 12'h666;
      20'h06a1e: out <= 12'h222;
      20'h06a1f: out <= 12'h666;
      20'h06a20: out <= 12'h222;
      20'h06a21: out <= 12'h666;
      20'h06a22: out <= 12'h222;
      20'h06a23: out <= 12'h666;
      20'h06a24: out <= 12'h222;
      20'h06a25: out <= 12'h222;
      20'h06a26: out <= 12'h222;
      20'h06a27: out <= 12'h222;
      20'h06a28: out <= 12'h000;
      20'h06a29: out <= 12'h000;
      20'h06a2a: out <= 12'h000;
      20'h06a2b: out <= 12'h666;
      20'h06a2c: out <= 12'h000;
      20'h06a2d: out <= 12'h666;
      20'h06a2e: out <= 12'h000;
      20'h06a2f: out <= 12'h666;
      20'h06a30: out <= 12'h000;
      20'h06a31: out <= 12'h666;
      20'h06a32: out <= 12'h000;
      20'h06a33: out <= 12'h666;
      20'h06a34: out <= 12'h000;
      20'h06a35: out <= 12'h000;
      20'h06a36: out <= 12'h000;
      20'h06a37: out <= 12'h000;
      20'h06a38: out <= 12'h222;
      20'h06a39: out <= 12'h222;
      20'h06a3a: out <= 12'h222;
      20'h06a3b: out <= 12'h222;
      20'h06a3c: out <= 12'h222;
      20'h06a3d: out <= 12'h222;
      20'h06a3e: out <= 12'h666;
      20'h06a3f: out <= 12'hbbb;
      20'h06a40: out <= 12'hfff;
      20'h06a41: out <= 12'hbbb;
      20'h06a42: out <= 12'h666;
      20'h06a43: out <= 12'h222;
      20'h06a44: out <= 12'h222;
      20'h06a45: out <= 12'h222;
      20'h06a46: out <= 12'h222;
      20'h06a47: out <= 12'h222;
      20'h06a48: out <= 12'h000;
      20'h06a49: out <= 12'h000;
      20'h06a4a: out <= 12'h000;
      20'h06a4b: out <= 12'h000;
      20'h06a4c: out <= 12'h000;
      20'h06a4d: out <= 12'h000;
      20'h06a4e: out <= 12'h666;
      20'h06a4f: out <= 12'hbbb;
      20'h06a50: out <= 12'hfff;
      20'h06a51: out <= 12'hbbb;
      20'h06a52: out <= 12'h666;
      20'h06a53: out <= 12'h000;
      20'h06a54: out <= 12'h000;
      20'h06a55: out <= 12'h000;
      20'h06a56: out <= 12'h000;
      20'h06a57: out <= 12'h000;
      20'h06a58: out <= 12'h222;
      20'h06a59: out <= 12'h222;
      20'h06a5a: out <= 12'h222;
      20'h06a5b: out <= 12'h222;
      20'h06a5c: out <= 12'h666;
      20'h06a5d: out <= 12'h222;
      20'h06a5e: out <= 12'h666;
      20'h06a5f: out <= 12'h222;
      20'h06a60: out <= 12'h666;
      20'h06a61: out <= 12'h222;
      20'h06a62: out <= 12'h666;
      20'h06a63: out <= 12'h222;
      20'h06a64: out <= 12'h666;
      20'h06a65: out <= 12'h222;
      20'h06a66: out <= 12'h222;
      20'h06a67: out <= 12'h222;
      20'h06a68: out <= 12'h000;
      20'h06a69: out <= 12'h000;
      20'h06a6a: out <= 12'h000;
      20'h06a6b: out <= 12'h000;
      20'h06a6c: out <= 12'h666;
      20'h06a6d: out <= 12'h000;
      20'h06a6e: out <= 12'h666;
      20'h06a6f: out <= 12'h000;
      20'h06a70: out <= 12'h666;
      20'h06a71: out <= 12'h000;
      20'h06a72: out <= 12'h666;
      20'h06a73: out <= 12'h000;
      20'h06a74: out <= 12'h666;
      20'h06a75: out <= 12'h000;
      20'h06a76: out <= 12'h000;
      20'h06a77: out <= 12'h000;
      20'h06a78: out <= 12'h222;
      20'h06a79: out <= 12'h222;
      20'h06a7a: out <= 12'h222;
      20'h06a7b: out <= 12'h222;
      20'h06a7c: out <= 12'h222;
      20'h06a7d: out <= 12'h222;
      20'h06a7e: out <= 12'h666;
      20'h06a7f: out <= 12'h666;
      20'h06a80: out <= 12'h666;
      20'h06a81: out <= 12'h666;
      20'h06a82: out <= 12'h666;
      20'h06a83: out <= 12'h222;
      20'h06a84: out <= 12'h222;
      20'h06a85: out <= 12'h222;
      20'h06a86: out <= 12'h222;
      20'h06a87: out <= 12'h222;
      20'h06a88: out <= 12'h000;
      20'h06a89: out <= 12'h000;
      20'h06a8a: out <= 12'h000;
      20'h06a8b: out <= 12'h000;
      20'h06a8c: out <= 12'h000;
      20'h06a8d: out <= 12'h000;
      20'h06a8e: out <= 12'h666;
      20'h06a8f: out <= 12'h666;
      20'h06a90: out <= 12'h666;
      20'h06a91: out <= 12'h666;
      20'h06a92: out <= 12'h666;
      20'h06a93: out <= 12'h000;
      20'h06a94: out <= 12'h000;
      20'h06a95: out <= 12'h000;
      20'h06a96: out <= 12'h000;
      20'h06a97: out <= 12'h000;
      20'h06a98: out <= 12'h603;
      20'h06a99: out <= 12'h603;
      20'h06a9a: out <= 12'h603;
      20'h06a9b: out <= 12'h603;
      20'h06a9c: out <= 12'h603;
      20'h06a9d: out <= 12'h603;
      20'h06a9e: out <= 12'h603;
      20'h06a9f: out <= 12'h603;
      20'h06aa0: out <= 12'h603;
      20'h06aa1: out <= 12'h603;
      20'h06aa2: out <= 12'h603;
      20'h06aa3: out <= 12'h603;
      20'h06aa4: out <= 12'hee9;
      20'h06aa5: out <= 12'hf87;
      20'h06aa6: out <= 12'hf87;
      20'h06aa7: out <= 12'hf87;
      20'h06aa8: out <= 12'hf87;
      20'h06aa9: out <= 12'hf87;
      20'h06aaa: out <= 12'hf87;
      20'h06aab: out <= 12'hb27;
      20'h06aac: out <= 12'hee9;
      20'h06aad: out <= 12'hf87;
      20'h06aae: out <= 12'hf87;
      20'h06aaf: out <= 12'hf87;
      20'h06ab0: out <= 12'hf87;
      20'h06ab1: out <= 12'hf87;
      20'h06ab2: out <= 12'hf87;
      20'h06ab3: out <= 12'hb27;
      20'h06ab4: out <= 12'hee9;
      20'h06ab5: out <= 12'hf87;
      20'h06ab6: out <= 12'hf87;
      20'h06ab7: out <= 12'hf87;
      20'h06ab8: out <= 12'hf87;
      20'h06ab9: out <= 12'hf87;
      20'h06aba: out <= 12'hf87;
      20'h06abb: out <= 12'hb27;
      20'h06abc: out <= 12'hee9;
      20'h06abd: out <= 12'hf87;
      20'h06abe: out <= 12'hf87;
      20'h06abf: out <= 12'hf87;
      20'h06ac0: out <= 12'hf87;
      20'h06ac1: out <= 12'hf87;
      20'h06ac2: out <= 12'hf87;
      20'h06ac3: out <= 12'hb27;
      20'h06ac4: out <= 12'h603;
      20'h06ac5: out <= 12'h603;
      20'h06ac6: out <= 12'h603;
      20'h06ac7: out <= 12'h603;
      20'h06ac8: out <= 12'h603;
      20'h06ac9: out <= 12'h603;
      20'h06aca: out <= 12'h603;
      20'h06acb: out <= 12'h603;
      20'h06acc: out <= 12'h603;
      20'h06acd: out <= 12'h603;
      20'h06ace: out <= 12'h603;
      20'h06acf: out <= 12'h603;
      20'h06ad0: out <= 12'h603;
      20'h06ad1: out <= 12'h603;
      20'h06ad2: out <= 12'h603;
      20'h06ad3: out <= 12'h603;
      20'h06ad4: out <= 12'h603;
      20'h06ad5: out <= 12'h603;
      20'h06ad6: out <= 12'h603;
      20'h06ad7: out <= 12'h603;
      20'h06ad8: out <= 12'h603;
      20'h06ad9: out <= 12'h603;
      20'h06ada: out <= 12'h603;
      20'h06adb: out <= 12'h603;
      20'h06adc: out <= 12'h603;
      20'h06add: out <= 12'h603;
      20'h06ade: out <= 12'h603;
      20'h06adf: out <= 12'h603;
      20'h06ae0: out <= 12'h603;
      20'h06ae1: out <= 12'h603;
      20'h06ae2: out <= 12'h603;
      20'h06ae3: out <= 12'h603;
      20'h06ae4: out <= 12'h603;
      20'h06ae5: out <= 12'h603;
      20'h06ae6: out <= 12'h603;
      20'h06ae7: out <= 12'h603;
      20'h06ae8: out <= 12'h603;
      20'h06ae9: out <= 12'h603;
      20'h06aea: out <= 12'h603;
      20'h06aeb: out <= 12'h603;
      20'h06aec: out <= 12'h603;
      20'h06aed: out <= 12'h603;
      20'h06aee: out <= 12'h603;
      20'h06aef: out <= 12'h603;
      20'h06af0: out <= 12'hee9;
      20'h06af1: out <= 12'hf87;
      20'h06af2: out <= 12'hf87;
      20'h06af3: out <= 12'hf87;
      20'h06af4: out <= 12'hf87;
      20'h06af5: out <= 12'hf87;
      20'h06af6: out <= 12'hf87;
      20'h06af7: out <= 12'hb27;
      20'h06af8: out <= 12'h000;
      20'h06af9: out <= 12'h000;
      20'h06afa: out <= 12'h000;
      20'h06afb: out <= 12'h000;
      20'h06afc: out <= 12'h000;
      20'h06afd: out <= 12'h000;
      20'h06afe: out <= 12'h000;
      20'h06aff: out <= 12'h000;
      20'h06b00: out <= 12'h777;
      20'h06b01: out <= 12'h777;
      20'h06b02: out <= 12'h555;
      20'h06b03: out <= 12'h555;
      20'h06b04: out <= 12'h555;
      20'h06b05: out <= 12'h555;
      20'h06b06: out <= 12'h555;
      20'h06b07: out <= 12'h555;
      20'h06b08: out <= 12'h555;
      20'h06b09: out <= 12'h555;
      20'h06b0a: out <= 12'h555;
      20'h06b0b: out <= 12'h555;
      20'h06b0c: out <= 12'h555;
      20'h06b0d: out <= 12'h555;
      20'h06b0e: out <= 12'h777;
      20'h06b0f: out <= 12'h777;
      20'h06b10: out <= 12'h000;
      20'h06b11: out <= 12'h000;
      20'h06b12: out <= 12'h000;
      20'h06b13: out <= 12'h000;
      20'h06b14: out <= 12'h000;
      20'h06b15: out <= 12'h000;
      20'h06b16: out <= 12'h000;
      20'h06b17: out <= 12'h000;
      20'h06b18: out <= 12'h000;
      20'h06b19: out <= 12'h000;
      20'h06b1a: out <= 12'h000;
      20'h06b1b: out <= 12'h000;
      20'h06b1c: out <= 12'h000;
      20'h06b1d: out <= 12'h000;
      20'h06b1e: out <= 12'h000;
      20'h06b1f: out <= 12'h000;
      20'h06b20: out <= 12'h000;
      20'h06b21: out <= 12'h000;
      20'h06b22: out <= 12'h000;
      20'h06b23: out <= 12'h000;
      20'h06b24: out <= 12'h000;
      20'h06b25: out <= 12'h000;
      20'h06b26: out <= 12'h000;
      20'h06b27: out <= 12'h000;
      20'h06b28: out <= 12'h000;
      20'h06b29: out <= 12'h000;
      20'h06b2a: out <= 12'h000;
      20'h06b2b: out <= 12'h000;
      20'h06b2c: out <= 12'h000;
      20'h06b2d: out <= 12'h000;
      20'h06b2e: out <= 12'h000;
      20'h06b2f: out <= 12'h000;
      20'h06b30: out <= 12'h222;
      20'h06b31: out <= 12'h222;
      20'h06b32: out <= 12'hbbb;
      20'h06b33: out <= 12'h666;
      20'h06b34: out <= 12'hbbb;
      20'h06b35: out <= 12'h666;
      20'h06b36: out <= 12'hbbb;
      20'h06b37: out <= 12'h666;
      20'h06b38: out <= 12'hbbb;
      20'h06b39: out <= 12'h666;
      20'h06b3a: out <= 12'hbbb;
      20'h06b3b: out <= 12'h666;
      20'h06b3c: out <= 12'hbbb;
      20'h06b3d: out <= 12'h222;
      20'h06b3e: out <= 12'h222;
      20'h06b3f: out <= 12'h222;
      20'h06b40: out <= 12'h000;
      20'h06b41: out <= 12'h000;
      20'h06b42: out <= 12'h666;
      20'h06b43: out <= 12'hbbb;
      20'h06b44: out <= 12'h666;
      20'h06b45: out <= 12'hbbb;
      20'h06b46: out <= 12'h666;
      20'h06b47: out <= 12'hbbb;
      20'h06b48: out <= 12'h666;
      20'h06b49: out <= 12'hbbb;
      20'h06b4a: out <= 12'h666;
      20'h06b4b: out <= 12'hbbb;
      20'h06b4c: out <= 12'h666;
      20'h06b4d: out <= 12'h000;
      20'h06b4e: out <= 12'h000;
      20'h06b4f: out <= 12'h000;
      20'h06b50: out <= 12'h222;
      20'h06b51: out <= 12'h222;
      20'h06b52: out <= 12'h222;
      20'h06b53: out <= 12'h222;
      20'h06b54: out <= 12'h222;
      20'h06b55: out <= 12'h222;
      20'h06b56: out <= 12'h666;
      20'h06b57: out <= 12'hbbb;
      20'h06b58: out <= 12'hfff;
      20'h06b59: out <= 12'hbbb;
      20'h06b5a: out <= 12'h666;
      20'h06b5b: out <= 12'h222;
      20'h06b5c: out <= 12'h222;
      20'h06b5d: out <= 12'h222;
      20'h06b5e: out <= 12'h222;
      20'h06b5f: out <= 12'h222;
      20'h06b60: out <= 12'h000;
      20'h06b61: out <= 12'h000;
      20'h06b62: out <= 12'h000;
      20'h06b63: out <= 12'h000;
      20'h06b64: out <= 12'h000;
      20'h06b65: out <= 12'h000;
      20'h06b66: out <= 12'h666;
      20'h06b67: out <= 12'hbbb;
      20'h06b68: out <= 12'hfff;
      20'h06b69: out <= 12'hbbb;
      20'h06b6a: out <= 12'h666;
      20'h06b6b: out <= 12'h000;
      20'h06b6c: out <= 12'h000;
      20'h06b6d: out <= 12'h000;
      20'h06b6e: out <= 12'h000;
      20'h06b6f: out <= 12'h000;
      20'h06b70: out <= 12'h222;
      20'h06b71: out <= 12'h222;
      20'h06b72: out <= 12'h222;
      20'h06b73: out <= 12'hbbb;
      20'h06b74: out <= 12'h666;
      20'h06b75: out <= 12'hbbb;
      20'h06b76: out <= 12'h666;
      20'h06b77: out <= 12'hbbb;
      20'h06b78: out <= 12'h666;
      20'h06b79: out <= 12'hbbb;
      20'h06b7a: out <= 12'h666;
      20'h06b7b: out <= 12'hbbb;
      20'h06b7c: out <= 12'h666;
      20'h06b7d: out <= 12'hbbb;
      20'h06b7e: out <= 12'h222;
      20'h06b7f: out <= 12'h222;
      20'h06b80: out <= 12'h000;
      20'h06b81: out <= 12'h000;
      20'h06b82: out <= 12'h000;
      20'h06b83: out <= 12'h666;
      20'h06b84: out <= 12'hbbb;
      20'h06b85: out <= 12'h666;
      20'h06b86: out <= 12'hbbb;
      20'h06b87: out <= 12'h666;
      20'h06b88: out <= 12'hbbb;
      20'h06b89: out <= 12'h666;
      20'h06b8a: out <= 12'hbbb;
      20'h06b8b: out <= 12'h666;
      20'h06b8c: out <= 12'hbbb;
      20'h06b8d: out <= 12'h666;
      20'h06b8e: out <= 12'h000;
      20'h06b8f: out <= 12'h000;
      20'h06b90: out <= 12'h222;
      20'h06b91: out <= 12'h222;
      20'h06b92: out <= 12'h222;
      20'h06b93: out <= 12'hbbb;
      20'h06b94: out <= 12'h222;
      20'h06b95: out <= 12'h666;
      20'h06b96: out <= 12'hfff;
      20'h06b97: out <= 12'hbbb;
      20'h06b98: out <= 12'hbbb;
      20'h06b99: out <= 12'hbbb;
      20'h06b9a: out <= 12'h666;
      20'h06b9b: out <= 12'h666;
      20'h06b9c: out <= 12'h222;
      20'h06b9d: out <= 12'hbbb;
      20'h06b9e: out <= 12'h222;
      20'h06b9f: out <= 12'h222;
      20'h06ba0: out <= 12'h000;
      20'h06ba1: out <= 12'h000;
      20'h06ba2: out <= 12'h000;
      20'h06ba3: out <= 12'h666;
      20'h06ba4: out <= 12'h000;
      20'h06ba5: out <= 12'h666;
      20'h06ba6: out <= 12'hfff;
      20'h06ba7: out <= 12'hbbb;
      20'h06ba8: out <= 12'hbbb;
      20'h06ba9: out <= 12'hbbb;
      20'h06baa: out <= 12'h666;
      20'h06bab: out <= 12'h666;
      20'h06bac: out <= 12'h000;
      20'h06bad: out <= 12'h666;
      20'h06bae: out <= 12'h000;
      20'h06baf: out <= 12'h000;
      20'h06bb0: out <= 12'h603;
      20'h06bb1: out <= 12'h603;
      20'h06bb2: out <= 12'h603;
      20'h06bb3: out <= 12'h603;
      20'h06bb4: out <= 12'h603;
      20'h06bb5: out <= 12'h603;
      20'h06bb6: out <= 12'h603;
      20'h06bb7: out <= 12'h603;
      20'h06bb8: out <= 12'h603;
      20'h06bb9: out <= 12'h603;
      20'h06bba: out <= 12'h603;
      20'h06bbb: out <= 12'h603;
      20'h06bbc: out <= 12'hee9;
      20'h06bbd: out <= 12'hf87;
      20'h06bbe: out <= 12'hee9;
      20'h06bbf: out <= 12'hee9;
      20'h06bc0: out <= 12'hee9;
      20'h06bc1: out <= 12'hb27;
      20'h06bc2: out <= 12'hf87;
      20'h06bc3: out <= 12'hb27;
      20'h06bc4: out <= 12'hee9;
      20'h06bc5: out <= 12'hf87;
      20'h06bc6: out <= 12'hee9;
      20'h06bc7: out <= 12'hee9;
      20'h06bc8: out <= 12'hee9;
      20'h06bc9: out <= 12'hb27;
      20'h06bca: out <= 12'hf87;
      20'h06bcb: out <= 12'hb27;
      20'h06bcc: out <= 12'hee9;
      20'h06bcd: out <= 12'hf87;
      20'h06bce: out <= 12'hee9;
      20'h06bcf: out <= 12'hee9;
      20'h06bd0: out <= 12'hee9;
      20'h06bd1: out <= 12'hb27;
      20'h06bd2: out <= 12'hf87;
      20'h06bd3: out <= 12'hb27;
      20'h06bd4: out <= 12'hee9;
      20'h06bd5: out <= 12'hf87;
      20'h06bd6: out <= 12'hee9;
      20'h06bd7: out <= 12'hee9;
      20'h06bd8: out <= 12'hee9;
      20'h06bd9: out <= 12'hb27;
      20'h06bda: out <= 12'hf87;
      20'h06bdb: out <= 12'hb27;
      20'h06bdc: out <= 12'h603;
      20'h06bdd: out <= 12'h603;
      20'h06bde: out <= 12'h603;
      20'h06bdf: out <= 12'h603;
      20'h06be0: out <= 12'h603;
      20'h06be1: out <= 12'h603;
      20'h06be2: out <= 12'h603;
      20'h06be3: out <= 12'h603;
      20'h06be4: out <= 12'h603;
      20'h06be5: out <= 12'h603;
      20'h06be6: out <= 12'h603;
      20'h06be7: out <= 12'h603;
      20'h06be8: out <= 12'h603;
      20'h06be9: out <= 12'h603;
      20'h06bea: out <= 12'h603;
      20'h06beb: out <= 12'h603;
      20'h06bec: out <= 12'h603;
      20'h06bed: out <= 12'h603;
      20'h06bee: out <= 12'h603;
      20'h06bef: out <= 12'h603;
      20'h06bf0: out <= 12'h603;
      20'h06bf1: out <= 12'h603;
      20'h06bf2: out <= 12'h603;
      20'h06bf3: out <= 12'h603;
      20'h06bf4: out <= 12'h603;
      20'h06bf5: out <= 12'h603;
      20'h06bf6: out <= 12'h603;
      20'h06bf7: out <= 12'h603;
      20'h06bf8: out <= 12'h603;
      20'h06bf9: out <= 12'h603;
      20'h06bfa: out <= 12'h603;
      20'h06bfb: out <= 12'h603;
      20'h06bfc: out <= 12'h603;
      20'h06bfd: out <= 12'h603;
      20'h06bfe: out <= 12'h603;
      20'h06bff: out <= 12'h603;
      20'h06c00: out <= 12'h603;
      20'h06c01: out <= 12'h603;
      20'h06c02: out <= 12'h603;
      20'h06c03: out <= 12'h603;
      20'h06c04: out <= 12'h603;
      20'h06c05: out <= 12'h603;
      20'h06c06: out <= 12'h603;
      20'h06c07: out <= 12'h603;
      20'h06c08: out <= 12'hee9;
      20'h06c09: out <= 12'hf87;
      20'h06c0a: out <= 12'hee9;
      20'h06c0b: out <= 12'hee9;
      20'h06c0c: out <= 12'hee9;
      20'h06c0d: out <= 12'hb27;
      20'h06c0e: out <= 12'hf87;
      20'h06c0f: out <= 12'hb27;
      20'h06c10: out <= 12'h000;
      20'h06c11: out <= 12'h000;
      20'h06c12: out <= 12'h000;
      20'h06c13: out <= 12'h000;
      20'h06c14: out <= 12'h000;
      20'h06c15: out <= 12'h000;
      20'h06c16: out <= 12'h000;
      20'h06c17: out <= 12'h000;
      20'h06c18: out <= 12'h777;
      20'h06c19: out <= 12'h555;
      20'h06c1a: out <= 12'h555;
      20'h06c1b: out <= 12'h555;
      20'h06c1c: out <= 12'h555;
      20'h06c1d: out <= 12'h555;
      20'h06c1e: out <= 12'h555;
      20'h06c1f: out <= 12'h555;
      20'h06c20: out <= 12'h555;
      20'h06c21: out <= 12'h555;
      20'h06c22: out <= 12'h555;
      20'h06c23: out <= 12'h555;
      20'h06c24: out <= 12'h555;
      20'h06c25: out <= 12'h555;
      20'h06c26: out <= 12'h555;
      20'h06c27: out <= 12'h777;
      20'h06c28: out <= 12'h000;
      20'h06c29: out <= 12'h000;
      20'h06c2a: out <= 12'h000;
      20'h06c2b: out <= 12'h000;
      20'h06c2c: out <= 12'h000;
      20'h06c2d: out <= 12'h000;
      20'h06c2e: out <= 12'h000;
      20'h06c2f: out <= 12'h000;
      20'h06c30: out <= 12'h000;
      20'h06c31: out <= 12'h000;
      20'h06c32: out <= 12'h000;
      20'h06c33: out <= 12'h000;
      20'h06c34: out <= 12'h000;
      20'h06c35: out <= 12'h000;
      20'h06c36: out <= 12'h000;
      20'h06c37: out <= 12'h000;
      20'h06c38: out <= 12'h000;
      20'h06c39: out <= 12'h000;
      20'h06c3a: out <= 12'h000;
      20'h06c3b: out <= 12'h000;
      20'h06c3c: out <= 12'h000;
      20'h06c3d: out <= 12'h000;
      20'h06c3e: out <= 12'h000;
      20'h06c3f: out <= 12'h000;
      20'h06c40: out <= 12'h000;
      20'h06c41: out <= 12'h000;
      20'h06c42: out <= 12'h000;
      20'h06c43: out <= 12'h000;
      20'h06c44: out <= 12'h000;
      20'h06c45: out <= 12'h000;
      20'h06c46: out <= 12'h000;
      20'h06c47: out <= 12'h000;
      20'h06c48: out <= 12'h222;
      20'h06c49: out <= 12'h222;
      20'h06c4a: out <= 12'h222;
      20'h06c4b: out <= 12'h666;
      20'h06c4c: out <= 12'h666;
      20'h06c4d: out <= 12'h666;
      20'h06c4e: out <= 12'h666;
      20'h06c4f: out <= 12'h666;
      20'h06c50: out <= 12'h666;
      20'h06c51: out <= 12'h666;
      20'h06c52: out <= 12'h666;
      20'h06c53: out <= 12'h666;
      20'h06c54: out <= 12'h222;
      20'h06c55: out <= 12'h222;
      20'h06c56: out <= 12'h222;
      20'h06c57: out <= 12'h222;
      20'h06c58: out <= 12'h000;
      20'h06c59: out <= 12'h000;
      20'h06c5a: out <= 12'h000;
      20'h06c5b: out <= 12'h666;
      20'h06c5c: out <= 12'h666;
      20'h06c5d: out <= 12'h666;
      20'h06c5e: out <= 12'h666;
      20'h06c5f: out <= 12'h666;
      20'h06c60: out <= 12'h666;
      20'h06c61: out <= 12'h666;
      20'h06c62: out <= 12'h666;
      20'h06c63: out <= 12'h666;
      20'h06c64: out <= 12'h000;
      20'h06c65: out <= 12'h000;
      20'h06c66: out <= 12'h000;
      20'h06c67: out <= 12'h000;
      20'h06c68: out <= 12'h222;
      20'h06c69: out <= 12'h222;
      20'h06c6a: out <= 12'h222;
      20'h06c6b: out <= 12'hbbb;
      20'h06c6c: out <= 12'h222;
      20'h06c6d: out <= 12'h666;
      20'h06c6e: out <= 12'h666;
      20'h06c6f: out <= 12'hbbb;
      20'h06c70: out <= 12'hfff;
      20'h06c71: out <= 12'hbbb;
      20'h06c72: out <= 12'h666;
      20'h06c73: out <= 12'h666;
      20'h06c74: out <= 12'h222;
      20'h06c75: out <= 12'hbbb;
      20'h06c76: out <= 12'h222;
      20'h06c77: out <= 12'h222;
      20'h06c78: out <= 12'h000;
      20'h06c79: out <= 12'h000;
      20'h06c7a: out <= 12'h000;
      20'h06c7b: out <= 12'h666;
      20'h06c7c: out <= 12'h000;
      20'h06c7d: out <= 12'h666;
      20'h06c7e: out <= 12'h666;
      20'h06c7f: out <= 12'hbbb;
      20'h06c80: out <= 12'hfff;
      20'h06c81: out <= 12'hbbb;
      20'h06c82: out <= 12'h666;
      20'h06c83: out <= 12'h666;
      20'h06c84: out <= 12'h000;
      20'h06c85: out <= 12'h666;
      20'h06c86: out <= 12'h000;
      20'h06c87: out <= 12'h000;
      20'h06c88: out <= 12'h222;
      20'h06c89: out <= 12'h222;
      20'h06c8a: out <= 12'h222;
      20'h06c8b: out <= 12'h222;
      20'h06c8c: out <= 12'h666;
      20'h06c8d: out <= 12'h666;
      20'h06c8e: out <= 12'h666;
      20'h06c8f: out <= 12'h666;
      20'h06c90: out <= 12'h666;
      20'h06c91: out <= 12'h666;
      20'h06c92: out <= 12'h666;
      20'h06c93: out <= 12'h666;
      20'h06c94: out <= 12'h666;
      20'h06c95: out <= 12'h222;
      20'h06c96: out <= 12'h222;
      20'h06c97: out <= 12'h222;
      20'h06c98: out <= 12'h000;
      20'h06c99: out <= 12'h000;
      20'h06c9a: out <= 12'h000;
      20'h06c9b: out <= 12'h000;
      20'h06c9c: out <= 12'h666;
      20'h06c9d: out <= 12'h666;
      20'h06c9e: out <= 12'h666;
      20'h06c9f: out <= 12'h666;
      20'h06ca0: out <= 12'h666;
      20'h06ca1: out <= 12'h666;
      20'h06ca2: out <= 12'h666;
      20'h06ca3: out <= 12'h666;
      20'h06ca4: out <= 12'h666;
      20'h06ca5: out <= 12'h000;
      20'h06ca6: out <= 12'h000;
      20'h06ca7: out <= 12'h000;
      20'h06ca8: out <= 12'h222;
      20'h06ca9: out <= 12'h222;
      20'h06caa: out <= 12'h666;
      20'h06cab: out <= 12'h666;
      20'h06cac: out <= 12'h666;
      20'h06cad: out <= 12'hfff;
      20'h06cae: out <= 12'hfff;
      20'h06caf: out <= 12'hbbb;
      20'h06cb0: out <= 12'hbbb;
      20'h06cb1: out <= 12'hbbb;
      20'h06cb2: out <= 12'h666;
      20'h06cb3: out <= 12'h666;
      20'h06cb4: out <= 12'h666;
      20'h06cb5: out <= 12'h666;
      20'h06cb6: out <= 12'h666;
      20'h06cb7: out <= 12'h222;
      20'h06cb8: out <= 12'h000;
      20'h06cb9: out <= 12'h000;
      20'h06cba: out <= 12'h666;
      20'h06cbb: out <= 12'hbbb;
      20'h06cbc: out <= 12'h666;
      20'h06cbd: out <= 12'hfff;
      20'h06cbe: out <= 12'hfff;
      20'h06cbf: out <= 12'hbbb;
      20'h06cc0: out <= 12'hbbb;
      20'h06cc1: out <= 12'hbbb;
      20'h06cc2: out <= 12'h666;
      20'h06cc3: out <= 12'h666;
      20'h06cc4: out <= 12'h666;
      20'h06cc5: out <= 12'hbbb;
      20'h06cc6: out <= 12'h666;
      20'h06cc7: out <= 12'h000;
      20'h06cc8: out <= 12'h603;
      20'h06cc9: out <= 12'h603;
      20'h06cca: out <= 12'h603;
      20'h06ccb: out <= 12'h603;
      20'h06ccc: out <= 12'h603;
      20'h06ccd: out <= 12'h603;
      20'h06cce: out <= 12'h603;
      20'h06ccf: out <= 12'h603;
      20'h06cd0: out <= 12'h603;
      20'h06cd1: out <= 12'h603;
      20'h06cd2: out <= 12'h603;
      20'h06cd3: out <= 12'h603;
      20'h06cd4: out <= 12'hee9;
      20'h06cd5: out <= 12'hf87;
      20'h06cd6: out <= 12'hee9;
      20'h06cd7: out <= 12'hf87;
      20'h06cd8: out <= 12'hf87;
      20'h06cd9: out <= 12'hb27;
      20'h06cda: out <= 12'hf87;
      20'h06cdb: out <= 12'hb27;
      20'h06cdc: out <= 12'hee9;
      20'h06cdd: out <= 12'hf87;
      20'h06cde: out <= 12'hee9;
      20'h06cdf: out <= 12'hf87;
      20'h06ce0: out <= 12'hf87;
      20'h06ce1: out <= 12'hb27;
      20'h06ce2: out <= 12'hf87;
      20'h06ce3: out <= 12'hb27;
      20'h06ce4: out <= 12'hee9;
      20'h06ce5: out <= 12'hf87;
      20'h06ce6: out <= 12'hee9;
      20'h06ce7: out <= 12'hf87;
      20'h06ce8: out <= 12'hf87;
      20'h06ce9: out <= 12'hb27;
      20'h06cea: out <= 12'hf87;
      20'h06ceb: out <= 12'hb27;
      20'h06cec: out <= 12'hee9;
      20'h06ced: out <= 12'hf87;
      20'h06cee: out <= 12'hee9;
      20'h06cef: out <= 12'hf87;
      20'h06cf0: out <= 12'hf87;
      20'h06cf1: out <= 12'hb27;
      20'h06cf2: out <= 12'hf87;
      20'h06cf3: out <= 12'hb27;
      20'h06cf4: out <= 12'h603;
      20'h06cf5: out <= 12'h603;
      20'h06cf6: out <= 12'h603;
      20'h06cf7: out <= 12'h603;
      20'h06cf8: out <= 12'h603;
      20'h06cf9: out <= 12'h603;
      20'h06cfa: out <= 12'h603;
      20'h06cfb: out <= 12'h603;
      20'h06cfc: out <= 12'h603;
      20'h06cfd: out <= 12'h603;
      20'h06cfe: out <= 12'h603;
      20'h06cff: out <= 12'h603;
      20'h06d00: out <= 12'h603;
      20'h06d01: out <= 12'h603;
      20'h06d02: out <= 12'h603;
      20'h06d03: out <= 12'h603;
      20'h06d04: out <= 12'h603;
      20'h06d05: out <= 12'h603;
      20'h06d06: out <= 12'h603;
      20'h06d07: out <= 12'h603;
      20'h06d08: out <= 12'h603;
      20'h06d09: out <= 12'h603;
      20'h06d0a: out <= 12'h603;
      20'h06d0b: out <= 12'h603;
      20'h06d0c: out <= 12'h603;
      20'h06d0d: out <= 12'h603;
      20'h06d0e: out <= 12'h603;
      20'h06d0f: out <= 12'h603;
      20'h06d10: out <= 12'h603;
      20'h06d11: out <= 12'h603;
      20'h06d12: out <= 12'h603;
      20'h06d13: out <= 12'h603;
      20'h06d14: out <= 12'h603;
      20'h06d15: out <= 12'h603;
      20'h06d16: out <= 12'h603;
      20'h06d17: out <= 12'h603;
      20'h06d18: out <= 12'h603;
      20'h06d19: out <= 12'h603;
      20'h06d1a: out <= 12'h603;
      20'h06d1b: out <= 12'h603;
      20'h06d1c: out <= 12'h603;
      20'h06d1d: out <= 12'h603;
      20'h06d1e: out <= 12'h603;
      20'h06d1f: out <= 12'h603;
      20'h06d20: out <= 12'hee9;
      20'h06d21: out <= 12'hf87;
      20'h06d22: out <= 12'hee9;
      20'h06d23: out <= 12'hf87;
      20'h06d24: out <= 12'hf87;
      20'h06d25: out <= 12'hb27;
      20'h06d26: out <= 12'hf87;
      20'h06d27: out <= 12'hb27;
      20'h06d28: out <= 12'h000;
      20'h06d29: out <= 12'h000;
      20'h06d2a: out <= 12'h000;
      20'h06d2b: out <= 12'h000;
      20'h06d2c: out <= 12'h000;
      20'h06d2d: out <= 12'h000;
      20'h06d2e: out <= 12'h000;
      20'h06d2f: out <= 12'h000;
      20'h06d30: out <= 12'h777;
      20'h06d31: out <= 12'h555;
      20'h06d32: out <= 12'h555;
      20'h06d33: out <= 12'h555;
      20'h06d34: out <= 12'h555;
      20'h06d35: out <= 12'h555;
      20'h06d36: out <= 12'h555;
      20'h06d37: out <= 12'h555;
      20'h06d38: out <= 12'h555;
      20'h06d39: out <= 12'h555;
      20'h06d3a: out <= 12'h555;
      20'h06d3b: out <= 12'h555;
      20'h06d3c: out <= 12'h555;
      20'h06d3d: out <= 12'h555;
      20'h06d3e: out <= 12'h555;
      20'h06d3f: out <= 12'h777;
      20'h06d40: out <= 12'h000;
      20'h06d41: out <= 12'h000;
      20'h06d42: out <= 12'h000;
      20'h06d43: out <= 12'h000;
      20'h06d44: out <= 12'h000;
      20'h06d45: out <= 12'h000;
      20'h06d46: out <= 12'h000;
      20'h06d47: out <= 12'h000;
      20'h06d48: out <= 12'h000;
      20'h06d49: out <= 12'h000;
      20'h06d4a: out <= 12'h000;
      20'h06d4b: out <= 12'h000;
      20'h06d4c: out <= 12'h000;
      20'h06d4d: out <= 12'h000;
      20'h06d4e: out <= 12'h000;
      20'h06d4f: out <= 12'h000;
      20'h06d50: out <= 12'h000;
      20'h06d51: out <= 12'h000;
      20'h06d52: out <= 12'h000;
      20'h06d53: out <= 12'h000;
      20'h06d54: out <= 12'h000;
      20'h06d55: out <= 12'h000;
      20'h06d56: out <= 12'h000;
      20'h06d57: out <= 12'h000;
      20'h06d58: out <= 12'h000;
      20'h06d59: out <= 12'h000;
      20'h06d5a: out <= 12'h000;
      20'h06d5b: out <= 12'h000;
      20'h06d5c: out <= 12'h000;
      20'h06d5d: out <= 12'h000;
      20'h06d5e: out <= 12'h000;
      20'h06d5f: out <= 12'h000;
      20'h06d60: out <= 12'h222;
      20'h06d61: out <= 12'h222;
      20'h06d62: out <= 12'h666;
      20'h06d63: out <= 12'hfff;
      20'h06d64: out <= 12'hfff;
      20'h06d65: out <= 12'hfff;
      20'h06d66: out <= 12'hfff;
      20'h06d67: out <= 12'hfff;
      20'h06d68: out <= 12'hfff;
      20'h06d69: out <= 12'hfff;
      20'h06d6a: out <= 12'hfff;
      20'h06d6b: out <= 12'hfff;
      20'h06d6c: out <= 12'h666;
      20'h06d6d: out <= 12'h222;
      20'h06d6e: out <= 12'h222;
      20'h06d6f: out <= 12'h222;
      20'h06d70: out <= 12'h000;
      20'h06d71: out <= 12'h000;
      20'h06d72: out <= 12'h666;
      20'h06d73: out <= 12'hfff;
      20'h06d74: out <= 12'hfff;
      20'h06d75: out <= 12'hfff;
      20'h06d76: out <= 12'hfff;
      20'h06d77: out <= 12'hfff;
      20'h06d78: out <= 12'hfff;
      20'h06d79: out <= 12'hfff;
      20'h06d7a: out <= 12'hfff;
      20'h06d7b: out <= 12'hfff;
      20'h06d7c: out <= 12'h666;
      20'h06d7d: out <= 12'h000;
      20'h06d7e: out <= 12'h000;
      20'h06d7f: out <= 12'h000;
      20'h06d80: out <= 12'h222;
      20'h06d81: out <= 12'h222;
      20'h06d82: out <= 12'h666;
      20'h06d83: out <= 12'h666;
      20'h06d84: out <= 12'h666;
      20'h06d85: out <= 12'hfff;
      20'h06d86: out <= 12'h666;
      20'h06d87: out <= 12'hbbb;
      20'h06d88: out <= 12'hfff;
      20'h06d89: out <= 12'hbbb;
      20'h06d8a: out <= 12'h666;
      20'h06d8b: out <= 12'h666;
      20'h06d8c: out <= 12'h666;
      20'h06d8d: out <= 12'h666;
      20'h06d8e: out <= 12'h666;
      20'h06d8f: out <= 12'h222;
      20'h06d90: out <= 12'h000;
      20'h06d91: out <= 12'h000;
      20'h06d92: out <= 12'h666;
      20'h06d93: out <= 12'hbbb;
      20'h06d94: out <= 12'h666;
      20'h06d95: out <= 12'hfff;
      20'h06d96: out <= 12'h666;
      20'h06d97: out <= 12'hbbb;
      20'h06d98: out <= 12'hfff;
      20'h06d99: out <= 12'hbbb;
      20'h06d9a: out <= 12'h666;
      20'h06d9b: out <= 12'h666;
      20'h06d9c: out <= 12'h666;
      20'h06d9d: out <= 12'hbbb;
      20'h06d9e: out <= 12'h666;
      20'h06d9f: out <= 12'h000;
      20'h06da0: out <= 12'h222;
      20'h06da1: out <= 12'h222;
      20'h06da2: out <= 12'h222;
      20'h06da3: out <= 12'h666;
      20'h06da4: out <= 12'hfff;
      20'h06da5: out <= 12'hfff;
      20'h06da6: out <= 12'hfff;
      20'h06da7: out <= 12'hfff;
      20'h06da8: out <= 12'hfff;
      20'h06da9: out <= 12'hfff;
      20'h06daa: out <= 12'hfff;
      20'h06dab: out <= 12'hfff;
      20'h06dac: out <= 12'hfff;
      20'h06dad: out <= 12'h666;
      20'h06dae: out <= 12'h222;
      20'h06daf: out <= 12'h222;
      20'h06db0: out <= 12'h000;
      20'h06db1: out <= 12'h000;
      20'h06db2: out <= 12'h000;
      20'h06db3: out <= 12'h666;
      20'h06db4: out <= 12'hfff;
      20'h06db5: out <= 12'hfff;
      20'h06db6: out <= 12'hfff;
      20'h06db7: out <= 12'hfff;
      20'h06db8: out <= 12'hfff;
      20'h06db9: out <= 12'hfff;
      20'h06dba: out <= 12'hfff;
      20'h06dbb: out <= 12'hfff;
      20'h06dbc: out <= 12'hfff;
      20'h06dbd: out <= 12'h666;
      20'h06dbe: out <= 12'h000;
      20'h06dbf: out <= 12'h000;
      20'h06dc0: out <= 12'h222;
      20'h06dc1: out <= 12'h222;
      20'h06dc2: out <= 12'h222;
      20'h06dc3: out <= 12'hbbb;
      20'h06dc4: out <= 12'h666;
      20'h06dc5: out <= 12'hfff;
      20'h06dc6: out <= 12'hfff;
      20'h06dc7: out <= 12'h666;
      20'h06dc8: out <= 12'h666;
      20'h06dc9: out <= 12'h666;
      20'h06dca: out <= 12'h666;
      20'h06dcb: out <= 12'h666;
      20'h06dcc: out <= 12'h666;
      20'h06dcd: out <= 12'hbbb;
      20'h06dce: out <= 12'h222;
      20'h06dcf: out <= 12'h222;
      20'h06dd0: out <= 12'h000;
      20'h06dd1: out <= 12'h000;
      20'h06dd2: out <= 12'h000;
      20'h06dd3: out <= 12'h666;
      20'h06dd4: out <= 12'h666;
      20'h06dd5: out <= 12'hfff;
      20'h06dd6: out <= 12'hfff;
      20'h06dd7: out <= 12'h666;
      20'h06dd8: out <= 12'h666;
      20'h06dd9: out <= 12'h666;
      20'h06dda: out <= 12'h666;
      20'h06ddb: out <= 12'h666;
      20'h06ddc: out <= 12'h666;
      20'h06ddd: out <= 12'h666;
      20'h06dde: out <= 12'h000;
      20'h06ddf: out <= 12'h000;
      20'h06de0: out <= 12'h603;
      20'h06de1: out <= 12'h603;
      20'h06de2: out <= 12'h603;
      20'h06de3: out <= 12'h603;
      20'h06de4: out <= 12'h603;
      20'h06de5: out <= 12'h603;
      20'h06de6: out <= 12'h603;
      20'h06de7: out <= 12'h603;
      20'h06de8: out <= 12'h603;
      20'h06de9: out <= 12'h603;
      20'h06dea: out <= 12'h603;
      20'h06deb: out <= 12'h603;
      20'h06dec: out <= 12'hee9;
      20'h06ded: out <= 12'hf87;
      20'h06dee: out <= 12'hee9;
      20'h06def: out <= 12'hf87;
      20'h06df0: out <= 12'hf87;
      20'h06df1: out <= 12'hb27;
      20'h06df2: out <= 12'hf87;
      20'h06df3: out <= 12'hb27;
      20'h06df4: out <= 12'hee9;
      20'h06df5: out <= 12'hf87;
      20'h06df6: out <= 12'hee9;
      20'h06df7: out <= 12'hf87;
      20'h06df8: out <= 12'hf87;
      20'h06df9: out <= 12'hb27;
      20'h06dfa: out <= 12'hf87;
      20'h06dfb: out <= 12'hb27;
      20'h06dfc: out <= 12'hee9;
      20'h06dfd: out <= 12'hf87;
      20'h06dfe: out <= 12'hee9;
      20'h06dff: out <= 12'hf87;
      20'h06e00: out <= 12'hf87;
      20'h06e01: out <= 12'hb27;
      20'h06e02: out <= 12'hf87;
      20'h06e03: out <= 12'hb27;
      20'h06e04: out <= 12'hee9;
      20'h06e05: out <= 12'hf87;
      20'h06e06: out <= 12'hee9;
      20'h06e07: out <= 12'hf87;
      20'h06e08: out <= 12'hf87;
      20'h06e09: out <= 12'hb27;
      20'h06e0a: out <= 12'hf87;
      20'h06e0b: out <= 12'hb27;
      20'h06e0c: out <= 12'h603;
      20'h06e0d: out <= 12'h603;
      20'h06e0e: out <= 12'h603;
      20'h06e0f: out <= 12'h603;
      20'h06e10: out <= 12'h603;
      20'h06e11: out <= 12'h603;
      20'h06e12: out <= 12'h603;
      20'h06e13: out <= 12'h603;
      20'h06e14: out <= 12'h603;
      20'h06e15: out <= 12'h603;
      20'h06e16: out <= 12'h603;
      20'h06e17: out <= 12'h603;
      20'h06e18: out <= 12'h603;
      20'h06e19: out <= 12'h603;
      20'h06e1a: out <= 12'h603;
      20'h06e1b: out <= 12'h603;
      20'h06e1c: out <= 12'h603;
      20'h06e1d: out <= 12'h603;
      20'h06e1e: out <= 12'h603;
      20'h06e1f: out <= 12'h603;
      20'h06e20: out <= 12'h603;
      20'h06e21: out <= 12'h603;
      20'h06e22: out <= 12'h603;
      20'h06e23: out <= 12'h603;
      20'h06e24: out <= 12'h603;
      20'h06e25: out <= 12'h603;
      20'h06e26: out <= 12'h603;
      20'h06e27: out <= 12'h603;
      20'h06e28: out <= 12'h603;
      20'h06e29: out <= 12'h603;
      20'h06e2a: out <= 12'h603;
      20'h06e2b: out <= 12'h603;
      20'h06e2c: out <= 12'h603;
      20'h06e2d: out <= 12'h603;
      20'h06e2e: out <= 12'h603;
      20'h06e2f: out <= 12'h603;
      20'h06e30: out <= 12'h603;
      20'h06e31: out <= 12'h603;
      20'h06e32: out <= 12'h603;
      20'h06e33: out <= 12'h603;
      20'h06e34: out <= 12'h603;
      20'h06e35: out <= 12'h603;
      20'h06e36: out <= 12'h603;
      20'h06e37: out <= 12'h603;
      20'h06e38: out <= 12'hee9;
      20'h06e39: out <= 12'hf87;
      20'h06e3a: out <= 12'hee9;
      20'h06e3b: out <= 12'hf87;
      20'h06e3c: out <= 12'hf87;
      20'h06e3d: out <= 12'hb27;
      20'h06e3e: out <= 12'hf87;
      20'h06e3f: out <= 12'hb27;
      20'h06e40: out <= 12'h000;
      20'h06e41: out <= 12'h000;
      20'h06e42: out <= 12'h000;
      20'h06e43: out <= 12'h000;
      20'h06e44: out <= 12'h000;
      20'h06e45: out <= 12'h000;
      20'h06e46: out <= 12'h000;
      20'h06e47: out <= 12'h000;
      20'h06e48: out <= 12'h777;
      20'h06e49: out <= 12'h555;
      20'h06e4a: out <= 12'h555;
      20'h06e4b: out <= 12'h555;
      20'h06e4c: out <= 12'h555;
      20'h06e4d: out <= 12'h555;
      20'h06e4e: out <= 12'h555;
      20'h06e4f: out <= 12'h555;
      20'h06e50: out <= 12'h555;
      20'h06e51: out <= 12'h555;
      20'h06e52: out <= 12'h555;
      20'h06e53: out <= 12'h555;
      20'h06e54: out <= 12'h555;
      20'h06e55: out <= 12'h555;
      20'h06e56: out <= 12'h555;
      20'h06e57: out <= 12'h777;
      20'h06e58: out <= 12'h000;
      20'h06e59: out <= 12'h000;
      20'h06e5a: out <= 12'h000;
      20'h06e5b: out <= 12'h000;
      20'h06e5c: out <= 12'h000;
      20'h06e5d: out <= 12'h000;
      20'h06e5e: out <= 12'h000;
      20'h06e5f: out <= 12'h000;
      20'h06e60: out <= 12'h000;
      20'h06e61: out <= 12'h000;
      20'h06e62: out <= 12'h000;
      20'h06e63: out <= 12'h000;
      20'h06e64: out <= 12'h000;
      20'h06e65: out <= 12'h000;
      20'h06e66: out <= 12'h000;
      20'h06e67: out <= 12'h000;
      20'h06e68: out <= 12'h000;
      20'h06e69: out <= 12'h000;
      20'h06e6a: out <= 12'h000;
      20'h06e6b: out <= 12'h000;
      20'h06e6c: out <= 12'h000;
      20'h06e6d: out <= 12'h000;
      20'h06e6e: out <= 12'h000;
      20'h06e6f: out <= 12'h000;
      20'h06e70: out <= 12'h000;
      20'h06e71: out <= 12'h000;
      20'h06e72: out <= 12'h000;
      20'h06e73: out <= 12'h000;
      20'h06e74: out <= 12'h000;
      20'h06e75: out <= 12'h000;
      20'h06e76: out <= 12'h000;
      20'h06e77: out <= 12'h000;
      20'h06e78: out <= 12'h222;
      20'h06e79: out <= 12'h666;
      20'h06e7a: out <= 12'hfff;
      20'h06e7b: out <= 12'hfff;
      20'h06e7c: out <= 12'hfff;
      20'h06e7d: out <= 12'h666;
      20'h06e7e: out <= 12'h666;
      20'h06e7f: out <= 12'h666;
      20'h06e80: out <= 12'hbbb;
      20'h06e81: out <= 12'h666;
      20'h06e82: out <= 12'h666;
      20'h06e83: out <= 12'h666;
      20'h06e84: out <= 12'h666;
      20'h06e85: out <= 12'h666;
      20'h06e86: out <= 12'h666;
      20'h06e87: out <= 12'h666;
      20'h06e88: out <= 12'h000;
      20'h06e89: out <= 12'h666;
      20'h06e8a: out <= 12'hfff;
      20'h06e8b: out <= 12'hfff;
      20'h06e8c: out <= 12'hfff;
      20'h06e8d: out <= 12'h666;
      20'h06e8e: out <= 12'h666;
      20'h06e8f: out <= 12'h666;
      20'h06e90: out <= 12'hbbb;
      20'h06e91: out <= 12'h666;
      20'h06e92: out <= 12'h666;
      20'h06e93: out <= 12'h666;
      20'h06e94: out <= 12'h666;
      20'h06e95: out <= 12'h666;
      20'h06e96: out <= 12'h666;
      20'h06e97: out <= 12'h666;
      20'h06e98: out <= 12'h222;
      20'h06e99: out <= 12'h222;
      20'h06e9a: out <= 12'h222;
      20'h06e9b: out <= 12'hbbb;
      20'h06e9c: out <= 12'h666;
      20'h06e9d: out <= 12'hfff;
      20'h06e9e: out <= 12'h666;
      20'h06e9f: out <= 12'hbbb;
      20'h06ea0: out <= 12'hfff;
      20'h06ea1: out <= 12'hbbb;
      20'h06ea2: out <= 12'h666;
      20'h06ea3: out <= 12'h666;
      20'h06ea4: out <= 12'h666;
      20'h06ea5: out <= 12'hbbb;
      20'h06ea6: out <= 12'h222;
      20'h06ea7: out <= 12'h222;
      20'h06ea8: out <= 12'h000;
      20'h06ea9: out <= 12'h000;
      20'h06eaa: out <= 12'h000;
      20'h06eab: out <= 12'h666;
      20'h06eac: out <= 12'h666;
      20'h06ead: out <= 12'hfff;
      20'h06eae: out <= 12'h666;
      20'h06eaf: out <= 12'hbbb;
      20'h06eb0: out <= 12'hfff;
      20'h06eb1: out <= 12'hbbb;
      20'h06eb2: out <= 12'h666;
      20'h06eb3: out <= 12'h666;
      20'h06eb4: out <= 12'h666;
      20'h06eb5: out <= 12'h666;
      20'h06eb6: out <= 12'h000;
      20'h06eb7: out <= 12'h000;
      20'h06eb8: out <= 12'h666;
      20'h06eb9: out <= 12'h666;
      20'h06eba: out <= 12'h666;
      20'h06ebb: out <= 12'h666;
      20'h06ebc: out <= 12'h666;
      20'h06ebd: out <= 12'h666;
      20'h06ebe: out <= 12'h666;
      20'h06ebf: out <= 12'hbbb;
      20'h06ec0: out <= 12'h666;
      20'h06ec1: out <= 12'h666;
      20'h06ec2: out <= 12'h666;
      20'h06ec3: out <= 12'hfff;
      20'h06ec4: out <= 12'hfff;
      20'h06ec5: out <= 12'hfff;
      20'h06ec6: out <= 12'h666;
      20'h06ec7: out <= 12'h222;
      20'h06ec8: out <= 12'h666;
      20'h06ec9: out <= 12'h666;
      20'h06eca: out <= 12'h666;
      20'h06ecb: out <= 12'h666;
      20'h06ecc: out <= 12'h666;
      20'h06ecd: out <= 12'h666;
      20'h06ece: out <= 12'h666;
      20'h06ecf: out <= 12'hbbb;
      20'h06ed0: out <= 12'h666;
      20'h06ed1: out <= 12'h666;
      20'h06ed2: out <= 12'h666;
      20'h06ed3: out <= 12'hfff;
      20'h06ed4: out <= 12'hfff;
      20'h06ed5: out <= 12'hfff;
      20'h06ed6: out <= 12'h666;
      20'h06ed7: out <= 12'h000;
      20'h06ed8: out <= 12'h222;
      20'h06ed9: out <= 12'h222;
      20'h06eda: out <= 12'h666;
      20'h06edb: out <= 12'h666;
      20'h06edc: out <= 12'h666;
      20'h06edd: out <= 12'hfff;
      20'h06ede: out <= 12'h666;
      20'h06edf: out <= 12'hbbb;
      20'h06ee0: out <= 12'hbbb;
      20'h06ee1: out <= 12'h666;
      20'h06ee2: out <= 12'h666;
      20'h06ee3: out <= 12'h666;
      20'h06ee4: out <= 12'h666;
      20'h06ee5: out <= 12'h666;
      20'h06ee6: out <= 12'h666;
      20'h06ee7: out <= 12'h222;
      20'h06ee8: out <= 12'h000;
      20'h06ee9: out <= 12'h000;
      20'h06eea: out <= 12'h666;
      20'h06eeb: out <= 12'hbbb;
      20'h06eec: out <= 12'h666;
      20'h06eed: out <= 12'hfff;
      20'h06eee: out <= 12'h666;
      20'h06eef: out <= 12'hbbb;
      20'h06ef0: out <= 12'hbbb;
      20'h06ef1: out <= 12'h666;
      20'h06ef2: out <= 12'h666;
      20'h06ef3: out <= 12'h666;
      20'h06ef4: out <= 12'h666;
      20'h06ef5: out <= 12'hbbb;
      20'h06ef6: out <= 12'h666;
      20'h06ef7: out <= 12'h000;
      20'h06ef8: out <= 12'h603;
      20'h06ef9: out <= 12'h603;
      20'h06efa: out <= 12'h603;
      20'h06efb: out <= 12'h603;
      20'h06efc: out <= 12'h603;
      20'h06efd: out <= 12'h603;
      20'h06efe: out <= 12'h603;
      20'h06eff: out <= 12'h603;
      20'h06f00: out <= 12'h603;
      20'h06f01: out <= 12'h603;
      20'h06f02: out <= 12'h603;
      20'h06f03: out <= 12'h603;
      20'h06f04: out <= 12'hee9;
      20'h06f05: out <= 12'hf87;
      20'h06f06: out <= 12'hee9;
      20'h06f07: out <= 12'hb27;
      20'h06f08: out <= 12'hb27;
      20'h06f09: out <= 12'hb27;
      20'h06f0a: out <= 12'hf87;
      20'h06f0b: out <= 12'hb27;
      20'h06f0c: out <= 12'hee9;
      20'h06f0d: out <= 12'hf87;
      20'h06f0e: out <= 12'hee9;
      20'h06f0f: out <= 12'hb27;
      20'h06f10: out <= 12'hb27;
      20'h06f11: out <= 12'hb27;
      20'h06f12: out <= 12'hf87;
      20'h06f13: out <= 12'hb27;
      20'h06f14: out <= 12'hee9;
      20'h06f15: out <= 12'hf87;
      20'h06f16: out <= 12'hee9;
      20'h06f17: out <= 12'hb27;
      20'h06f18: out <= 12'hb27;
      20'h06f19: out <= 12'hb27;
      20'h06f1a: out <= 12'hf87;
      20'h06f1b: out <= 12'hb27;
      20'h06f1c: out <= 12'hee9;
      20'h06f1d: out <= 12'hf87;
      20'h06f1e: out <= 12'hee9;
      20'h06f1f: out <= 12'hb27;
      20'h06f20: out <= 12'hb27;
      20'h06f21: out <= 12'hb27;
      20'h06f22: out <= 12'hf87;
      20'h06f23: out <= 12'hb27;
      20'h06f24: out <= 12'h603;
      20'h06f25: out <= 12'h603;
      20'h06f26: out <= 12'h603;
      20'h06f27: out <= 12'h603;
      20'h06f28: out <= 12'h603;
      20'h06f29: out <= 12'h603;
      20'h06f2a: out <= 12'h603;
      20'h06f2b: out <= 12'h603;
      20'h06f2c: out <= 12'h603;
      20'h06f2d: out <= 12'h603;
      20'h06f2e: out <= 12'h603;
      20'h06f2f: out <= 12'h603;
      20'h06f30: out <= 12'h603;
      20'h06f31: out <= 12'h603;
      20'h06f32: out <= 12'h603;
      20'h06f33: out <= 12'h603;
      20'h06f34: out <= 12'h603;
      20'h06f35: out <= 12'h603;
      20'h06f36: out <= 12'h603;
      20'h06f37: out <= 12'h603;
      20'h06f38: out <= 12'h603;
      20'h06f39: out <= 12'h603;
      20'h06f3a: out <= 12'h603;
      20'h06f3b: out <= 12'h603;
      20'h06f3c: out <= 12'h603;
      20'h06f3d: out <= 12'h603;
      20'h06f3e: out <= 12'h603;
      20'h06f3f: out <= 12'h603;
      20'h06f40: out <= 12'h603;
      20'h06f41: out <= 12'h603;
      20'h06f42: out <= 12'h603;
      20'h06f43: out <= 12'h603;
      20'h06f44: out <= 12'h603;
      20'h06f45: out <= 12'h603;
      20'h06f46: out <= 12'h603;
      20'h06f47: out <= 12'h603;
      20'h06f48: out <= 12'h603;
      20'h06f49: out <= 12'h603;
      20'h06f4a: out <= 12'h603;
      20'h06f4b: out <= 12'h603;
      20'h06f4c: out <= 12'h603;
      20'h06f4d: out <= 12'h603;
      20'h06f4e: out <= 12'h603;
      20'h06f4f: out <= 12'h603;
      20'h06f50: out <= 12'hee9;
      20'h06f51: out <= 12'hf87;
      20'h06f52: out <= 12'hee9;
      20'h06f53: out <= 12'hb27;
      20'h06f54: out <= 12'hb27;
      20'h06f55: out <= 12'hb27;
      20'h06f56: out <= 12'hf87;
      20'h06f57: out <= 12'hb27;
      20'h06f58: out <= 12'h000;
      20'h06f59: out <= 12'h000;
      20'h06f5a: out <= 12'h000;
      20'h06f5b: out <= 12'h000;
      20'h06f5c: out <= 12'h000;
      20'h06f5d: out <= 12'h000;
      20'h06f5e: out <= 12'h000;
      20'h06f5f: out <= 12'h000;
      20'h06f60: out <= 12'h777;
      20'h06f61: out <= 12'h555;
      20'h06f62: out <= 12'h555;
      20'h06f63: out <= 12'h555;
      20'h06f64: out <= 12'h555;
      20'h06f65: out <= 12'h555;
      20'h06f66: out <= 12'h555;
      20'h06f67: out <= 12'h555;
      20'h06f68: out <= 12'h555;
      20'h06f69: out <= 12'h555;
      20'h06f6a: out <= 12'h555;
      20'h06f6b: out <= 12'h555;
      20'h06f6c: out <= 12'h555;
      20'h06f6d: out <= 12'h555;
      20'h06f6e: out <= 12'h555;
      20'h06f6f: out <= 12'h777;
      20'h06f70: out <= 12'h000;
      20'h06f71: out <= 12'h000;
      20'h06f72: out <= 12'h000;
      20'h06f73: out <= 12'h000;
      20'h06f74: out <= 12'h000;
      20'h06f75: out <= 12'h000;
      20'h06f76: out <= 12'h000;
      20'h06f77: out <= 12'h000;
      20'h06f78: out <= 12'h000;
      20'h06f79: out <= 12'h000;
      20'h06f7a: out <= 12'h000;
      20'h06f7b: out <= 12'h000;
      20'h06f7c: out <= 12'h000;
      20'h06f7d: out <= 12'h000;
      20'h06f7e: out <= 12'h000;
      20'h06f7f: out <= 12'h000;
      20'h06f80: out <= 12'h000;
      20'h06f81: out <= 12'h000;
      20'h06f82: out <= 12'h000;
      20'h06f83: out <= 12'h000;
      20'h06f84: out <= 12'h000;
      20'h06f85: out <= 12'h000;
      20'h06f86: out <= 12'h000;
      20'h06f87: out <= 12'h000;
      20'h06f88: out <= 12'h000;
      20'h06f89: out <= 12'h000;
      20'h06f8a: out <= 12'h000;
      20'h06f8b: out <= 12'h000;
      20'h06f8c: out <= 12'h000;
      20'h06f8d: out <= 12'h000;
      20'h06f8e: out <= 12'h000;
      20'h06f8f: out <= 12'h000;
      20'h06f90: out <= 12'h222;
      20'h06f91: out <= 12'h666;
      20'h06f92: out <= 12'hbbb;
      20'h06f93: out <= 12'hbbb;
      20'h06f94: out <= 12'h666;
      20'h06f95: out <= 12'hbbb;
      20'h06f96: out <= 12'hfff;
      20'h06f97: out <= 12'hfff;
      20'h06f98: out <= 12'h666;
      20'h06f99: out <= 12'hbbb;
      20'h06f9a: out <= 12'hbbb;
      20'h06f9b: out <= 12'hbbb;
      20'h06f9c: out <= 12'hbbb;
      20'h06f9d: out <= 12'hbbb;
      20'h06f9e: out <= 12'hbbb;
      20'h06f9f: out <= 12'hbbb;
      20'h06fa0: out <= 12'h000;
      20'h06fa1: out <= 12'h666;
      20'h06fa2: out <= 12'hbbb;
      20'h06fa3: out <= 12'hbbb;
      20'h06fa4: out <= 12'h666;
      20'h06fa5: out <= 12'hbbb;
      20'h06fa6: out <= 12'hfff;
      20'h06fa7: out <= 12'hfff;
      20'h06fa8: out <= 12'h666;
      20'h06fa9: out <= 12'hbbb;
      20'h06faa: out <= 12'hbbb;
      20'h06fab: out <= 12'hbbb;
      20'h06fac: out <= 12'hbbb;
      20'h06fad: out <= 12'hbbb;
      20'h06fae: out <= 12'hbbb;
      20'h06faf: out <= 12'hbbb;
      20'h06fb0: out <= 12'h222;
      20'h06fb1: out <= 12'h222;
      20'h06fb2: out <= 12'h666;
      20'h06fb3: out <= 12'h666;
      20'h06fb4: out <= 12'h666;
      20'h06fb5: out <= 12'hfff;
      20'h06fb6: out <= 12'h666;
      20'h06fb7: out <= 12'hbbb;
      20'h06fb8: out <= 12'hfff;
      20'h06fb9: out <= 12'hbbb;
      20'h06fba: out <= 12'h666;
      20'h06fbb: out <= 12'h666;
      20'h06fbc: out <= 12'h666;
      20'h06fbd: out <= 12'h666;
      20'h06fbe: out <= 12'h666;
      20'h06fbf: out <= 12'h222;
      20'h06fc0: out <= 12'h000;
      20'h06fc1: out <= 12'h000;
      20'h06fc2: out <= 12'h666;
      20'h06fc3: out <= 12'hbbb;
      20'h06fc4: out <= 12'h666;
      20'h06fc5: out <= 12'hfff;
      20'h06fc6: out <= 12'h666;
      20'h06fc7: out <= 12'hbbb;
      20'h06fc8: out <= 12'hfff;
      20'h06fc9: out <= 12'hbbb;
      20'h06fca: out <= 12'h666;
      20'h06fcb: out <= 12'h666;
      20'h06fcc: out <= 12'h666;
      20'h06fcd: out <= 12'hbbb;
      20'h06fce: out <= 12'h666;
      20'h06fcf: out <= 12'h000;
      20'h06fd0: out <= 12'hbbb;
      20'h06fd1: out <= 12'hbbb;
      20'h06fd2: out <= 12'hbbb;
      20'h06fd3: out <= 12'hbbb;
      20'h06fd4: out <= 12'hbbb;
      20'h06fd5: out <= 12'hbbb;
      20'h06fd6: out <= 12'hbbb;
      20'h06fd7: out <= 12'h666;
      20'h06fd8: out <= 12'hfff;
      20'h06fd9: out <= 12'hfff;
      20'h06fda: out <= 12'hbbb;
      20'h06fdb: out <= 12'h666;
      20'h06fdc: out <= 12'hbbb;
      20'h06fdd: out <= 12'hbbb;
      20'h06fde: out <= 12'h666;
      20'h06fdf: out <= 12'h222;
      20'h06fe0: out <= 12'hbbb;
      20'h06fe1: out <= 12'hbbb;
      20'h06fe2: out <= 12'hbbb;
      20'h06fe3: out <= 12'hbbb;
      20'h06fe4: out <= 12'hbbb;
      20'h06fe5: out <= 12'hbbb;
      20'h06fe6: out <= 12'hbbb;
      20'h06fe7: out <= 12'h666;
      20'h06fe8: out <= 12'hfff;
      20'h06fe9: out <= 12'hfff;
      20'h06fea: out <= 12'hbbb;
      20'h06feb: out <= 12'h666;
      20'h06fec: out <= 12'hbbb;
      20'h06fed: out <= 12'hbbb;
      20'h06fee: out <= 12'h666;
      20'h06fef: out <= 12'h000;
      20'h06ff0: out <= 12'h222;
      20'h06ff1: out <= 12'h222;
      20'h06ff2: out <= 12'h222;
      20'h06ff3: out <= 12'hbbb;
      20'h06ff4: out <= 12'h666;
      20'h06ff5: out <= 12'hfff;
      20'h06ff6: out <= 12'h666;
      20'h06ff7: out <= 12'hfff;
      20'h06ff8: out <= 12'hbbb;
      20'h06ff9: out <= 12'hbbb;
      20'h06ffa: out <= 12'h666;
      20'h06ffb: out <= 12'h666;
      20'h06ffc: out <= 12'h666;
      20'h06ffd: out <= 12'hbbb;
      20'h06ffe: out <= 12'h222;
      20'h06fff: out <= 12'h222;
      20'h07000: out <= 12'h000;
      20'h07001: out <= 12'h000;
      20'h07002: out <= 12'h000;
      20'h07003: out <= 12'h666;
      20'h07004: out <= 12'h666;
      20'h07005: out <= 12'hfff;
      20'h07006: out <= 12'h666;
      20'h07007: out <= 12'hfff;
      20'h07008: out <= 12'hbbb;
      20'h07009: out <= 12'hbbb;
      20'h0700a: out <= 12'h666;
      20'h0700b: out <= 12'h666;
      20'h0700c: out <= 12'h666;
      20'h0700d: out <= 12'h666;
      20'h0700e: out <= 12'h000;
      20'h0700f: out <= 12'h000;
      20'h07010: out <= 12'h603;
      20'h07011: out <= 12'h603;
      20'h07012: out <= 12'h603;
      20'h07013: out <= 12'h603;
      20'h07014: out <= 12'h603;
      20'h07015: out <= 12'h603;
      20'h07016: out <= 12'h603;
      20'h07017: out <= 12'h603;
      20'h07018: out <= 12'h603;
      20'h07019: out <= 12'h603;
      20'h0701a: out <= 12'h603;
      20'h0701b: out <= 12'h603;
      20'h0701c: out <= 12'hee9;
      20'h0701d: out <= 12'hf87;
      20'h0701e: out <= 12'hf87;
      20'h0701f: out <= 12'hf87;
      20'h07020: out <= 12'hf87;
      20'h07021: out <= 12'hf87;
      20'h07022: out <= 12'hf87;
      20'h07023: out <= 12'hb27;
      20'h07024: out <= 12'hee9;
      20'h07025: out <= 12'hf87;
      20'h07026: out <= 12'hf87;
      20'h07027: out <= 12'hf87;
      20'h07028: out <= 12'hf87;
      20'h07029: out <= 12'hf87;
      20'h0702a: out <= 12'hf87;
      20'h0702b: out <= 12'hb27;
      20'h0702c: out <= 12'hee9;
      20'h0702d: out <= 12'hf87;
      20'h0702e: out <= 12'hf87;
      20'h0702f: out <= 12'hf87;
      20'h07030: out <= 12'hf87;
      20'h07031: out <= 12'hf87;
      20'h07032: out <= 12'hf87;
      20'h07033: out <= 12'hb27;
      20'h07034: out <= 12'hee9;
      20'h07035: out <= 12'hf87;
      20'h07036: out <= 12'hf87;
      20'h07037: out <= 12'hf87;
      20'h07038: out <= 12'hf87;
      20'h07039: out <= 12'hf87;
      20'h0703a: out <= 12'hf87;
      20'h0703b: out <= 12'hb27;
      20'h0703c: out <= 12'h603;
      20'h0703d: out <= 12'h603;
      20'h0703e: out <= 12'h603;
      20'h0703f: out <= 12'h603;
      20'h07040: out <= 12'h603;
      20'h07041: out <= 12'h603;
      20'h07042: out <= 12'h603;
      20'h07043: out <= 12'h603;
      20'h07044: out <= 12'h603;
      20'h07045: out <= 12'h603;
      20'h07046: out <= 12'h603;
      20'h07047: out <= 12'h603;
      20'h07048: out <= 12'h603;
      20'h07049: out <= 12'h603;
      20'h0704a: out <= 12'h603;
      20'h0704b: out <= 12'h603;
      20'h0704c: out <= 12'h603;
      20'h0704d: out <= 12'h603;
      20'h0704e: out <= 12'h603;
      20'h0704f: out <= 12'h603;
      20'h07050: out <= 12'h603;
      20'h07051: out <= 12'h603;
      20'h07052: out <= 12'h603;
      20'h07053: out <= 12'h603;
      20'h07054: out <= 12'h603;
      20'h07055: out <= 12'h603;
      20'h07056: out <= 12'h603;
      20'h07057: out <= 12'h603;
      20'h07058: out <= 12'h603;
      20'h07059: out <= 12'h603;
      20'h0705a: out <= 12'h603;
      20'h0705b: out <= 12'h603;
      20'h0705c: out <= 12'h603;
      20'h0705d: out <= 12'h603;
      20'h0705e: out <= 12'h603;
      20'h0705f: out <= 12'h603;
      20'h07060: out <= 12'h603;
      20'h07061: out <= 12'h603;
      20'h07062: out <= 12'h603;
      20'h07063: out <= 12'h603;
      20'h07064: out <= 12'h603;
      20'h07065: out <= 12'h603;
      20'h07066: out <= 12'h603;
      20'h07067: out <= 12'h603;
      20'h07068: out <= 12'hee9;
      20'h07069: out <= 12'hf87;
      20'h0706a: out <= 12'hf87;
      20'h0706b: out <= 12'hf87;
      20'h0706c: out <= 12'hf87;
      20'h0706d: out <= 12'hf87;
      20'h0706e: out <= 12'hf87;
      20'h0706f: out <= 12'hb27;
      20'h07070: out <= 12'h000;
      20'h07071: out <= 12'h000;
      20'h07072: out <= 12'h000;
      20'h07073: out <= 12'h000;
      20'h07074: out <= 12'h000;
      20'h07075: out <= 12'h000;
      20'h07076: out <= 12'h000;
      20'h07077: out <= 12'h000;
      20'h07078: out <= 12'h777;
      20'h07079: out <= 12'h555;
      20'h0707a: out <= 12'h555;
      20'h0707b: out <= 12'h555;
      20'h0707c: out <= 12'h555;
      20'h0707d: out <= 12'h555;
      20'h0707e: out <= 12'h555;
      20'h0707f: out <= 12'h555;
      20'h07080: out <= 12'h555;
      20'h07081: out <= 12'h555;
      20'h07082: out <= 12'h555;
      20'h07083: out <= 12'h555;
      20'h07084: out <= 12'h555;
      20'h07085: out <= 12'h555;
      20'h07086: out <= 12'h555;
      20'h07087: out <= 12'h777;
      20'h07088: out <= 12'h000;
      20'h07089: out <= 12'h000;
      20'h0708a: out <= 12'h000;
      20'h0708b: out <= 12'h000;
      20'h0708c: out <= 12'h000;
      20'h0708d: out <= 12'h000;
      20'h0708e: out <= 12'h000;
      20'h0708f: out <= 12'h000;
      20'h07090: out <= 12'h000;
      20'h07091: out <= 12'h000;
      20'h07092: out <= 12'h000;
      20'h07093: out <= 12'h000;
      20'h07094: out <= 12'h000;
      20'h07095: out <= 12'h000;
      20'h07096: out <= 12'h000;
      20'h07097: out <= 12'h000;
      20'h07098: out <= 12'h000;
      20'h07099: out <= 12'h000;
      20'h0709a: out <= 12'h000;
      20'h0709b: out <= 12'h000;
      20'h0709c: out <= 12'h000;
      20'h0709d: out <= 12'h000;
      20'h0709e: out <= 12'h000;
      20'h0709f: out <= 12'h000;
      20'h070a0: out <= 12'h000;
      20'h070a1: out <= 12'h000;
      20'h070a2: out <= 12'h000;
      20'h070a3: out <= 12'h000;
      20'h070a4: out <= 12'h000;
      20'h070a5: out <= 12'h000;
      20'h070a6: out <= 12'h000;
      20'h070a7: out <= 12'h000;
      20'h070a8: out <= 12'h222;
      20'h070a9: out <= 12'h666;
      20'h070aa: out <= 12'hbbb;
      20'h070ab: out <= 12'hbbb;
      20'h070ac: out <= 12'h666;
      20'h070ad: out <= 12'hbbb;
      20'h070ae: out <= 12'hbbb;
      20'h070af: out <= 12'hfff;
      20'h070b0: out <= 12'h666;
      20'h070b1: out <= 12'hfff;
      20'h070b2: out <= 12'hfff;
      20'h070b3: out <= 12'hfff;
      20'h070b4: out <= 12'hfff;
      20'h070b5: out <= 12'hfff;
      20'h070b6: out <= 12'hfff;
      20'h070b7: out <= 12'hfff;
      20'h070b8: out <= 12'h000;
      20'h070b9: out <= 12'h666;
      20'h070ba: out <= 12'hbbb;
      20'h070bb: out <= 12'hbbb;
      20'h070bc: out <= 12'h666;
      20'h070bd: out <= 12'hbbb;
      20'h070be: out <= 12'hbbb;
      20'h070bf: out <= 12'hfff;
      20'h070c0: out <= 12'h666;
      20'h070c1: out <= 12'hfff;
      20'h070c2: out <= 12'hfff;
      20'h070c3: out <= 12'hfff;
      20'h070c4: out <= 12'hfff;
      20'h070c5: out <= 12'hfff;
      20'h070c6: out <= 12'hfff;
      20'h070c7: out <= 12'hfff;
      20'h070c8: out <= 12'h222;
      20'h070c9: out <= 12'h222;
      20'h070ca: out <= 12'h222;
      20'h070cb: out <= 12'hbbb;
      20'h070cc: out <= 12'h666;
      20'h070cd: out <= 12'hfff;
      20'h070ce: out <= 12'hbbb;
      20'h070cf: out <= 12'h666;
      20'h070d0: out <= 12'h666;
      20'h070d1: out <= 12'h666;
      20'h070d2: out <= 12'h666;
      20'h070d3: out <= 12'h666;
      20'h070d4: out <= 12'h666;
      20'h070d5: out <= 12'hbbb;
      20'h070d6: out <= 12'h222;
      20'h070d7: out <= 12'h222;
      20'h070d8: out <= 12'h000;
      20'h070d9: out <= 12'h000;
      20'h070da: out <= 12'h000;
      20'h070db: out <= 12'h666;
      20'h070dc: out <= 12'h666;
      20'h070dd: out <= 12'hfff;
      20'h070de: out <= 12'hbbb;
      20'h070df: out <= 12'h666;
      20'h070e0: out <= 12'h666;
      20'h070e1: out <= 12'h666;
      20'h070e2: out <= 12'h666;
      20'h070e3: out <= 12'h666;
      20'h070e4: out <= 12'h666;
      20'h070e5: out <= 12'h666;
      20'h070e6: out <= 12'h000;
      20'h070e7: out <= 12'h000;
      20'h070e8: out <= 12'hfff;
      20'h070e9: out <= 12'hfff;
      20'h070ea: out <= 12'hfff;
      20'h070eb: out <= 12'hfff;
      20'h070ec: out <= 12'hfff;
      20'h070ed: out <= 12'hfff;
      20'h070ee: out <= 12'hfff;
      20'h070ef: out <= 12'h666;
      20'h070f0: out <= 12'hfff;
      20'h070f1: out <= 12'hbbb;
      20'h070f2: out <= 12'hbbb;
      20'h070f3: out <= 12'h666;
      20'h070f4: out <= 12'hbbb;
      20'h070f5: out <= 12'hbbb;
      20'h070f6: out <= 12'h666;
      20'h070f7: out <= 12'h222;
      20'h070f8: out <= 12'hfff;
      20'h070f9: out <= 12'hfff;
      20'h070fa: out <= 12'hfff;
      20'h070fb: out <= 12'hfff;
      20'h070fc: out <= 12'hfff;
      20'h070fd: out <= 12'hfff;
      20'h070fe: out <= 12'hfff;
      20'h070ff: out <= 12'h666;
      20'h07100: out <= 12'hfff;
      20'h07101: out <= 12'hbbb;
      20'h07102: out <= 12'hbbb;
      20'h07103: out <= 12'h666;
      20'h07104: out <= 12'hbbb;
      20'h07105: out <= 12'hbbb;
      20'h07106: out <= 12'h666;
      20'h07107: out <= 12'h000;
      20'h07108: out <= 12'h222;
      20'h07109: out <= 12'h222;
      20'h0710a: out <= 12'h666;
      20'h0710b: out <= 12'h666;
      20'h0710c: out <= 12'h666;
      20'h0710d: out <= 12'hfff;
      20'h0710e: out <= 12'h666;
      20'h0710f: out <= 12'hfff;
      20'h07110: out <= 12'hfff;
      20'h07111: out <= 12'hbbb;
      20'h07112: out <= 12'h666;
      20'h07113: out <= 12'h666;
      20'h07114: out <= 12'h666;
      20'h07115: out <= 12'h666;
      20'h07116: out <= 12'h666;
      20'h07117: out <= 12'h222;
      20'h07118: out <= 12'h000;
      20'h07119: out <= 12'h000;
      20'h0711a: out <= 12'h666;
      20'h0711b: out <= 12'hbbb;
      20'h0711c: out <= 12'h666;
      20'h0711d: out <= 12'hfff;
      20'h0711e: out <= 12'h666;
      20'h0711f: out <= 12'hfff;
      20'h07120: out <= 12'hfff;
      20'h07121: out <= 12'hbbb;
      20'h07122: out <= 12'h666;
      20'h07123: out <= 12'h666;
      20'h07124: out <= 12'h666;
      20'h07125: out <= 12'hbbb;
      20'h07126: out <= 12'h666;
      20'h07127: out <= 12'h000;
      20'h07128: out <= 12'h603;
      20'h07129: out <= 12'h603;
      20'h0712a: out <= 12'h603;
      20'h0712b: out <= 12'h603;
      20'h0712c: out <= 12'h603;
      20'h0712d: out <= 12'h603;
      20'h0712e: out <= 12'h603;
      20'h0712f: out <= 12'h603;
      20'h07130: out <= 12'h603;
      20'h07131: out <= 12'h603;
      20'h07132: out <= 12'h603;
      20'h07133: out <= 12'h603;
      20'h07134: out <= 12'hb27;
      20'h07135: out <= 12'hb27;
      20'h07136: out <= 12'hb27;
      20'h07137: out <= 12'hb27;
      20'h07138: out <= 12'hb27;
      20'h07139: out <= 12'hb27;
      20'h0713a: out <= 12'hb27;
      20'h0713b: out <= 12'hb27;
      20'h0713c: out <= 12'hb27;
      20'h0713d: out <= 12'hb27;
      20'h0713e: out <= 12'hb27;
      20'h0713f: out <= 12'hb27;
      20'h07140: out <= 12'hb27;
      20'h07141: out <= 12'hb27;
      20'h07142: out <= 12'hb27;
      20'h07143: out <= 12'hb27;
      20'h07144: out <= 12'hb27;
      20'h07145: out <= 12'hb27;
      20'h07146: out <= 12'hb27;
      20'h07147: out <= 12'hb27;
      20'h07148: out <= 12'hb27;
      20'h07149: out <= 12'hb27;
      20'h0714a: out <= 12'hb27;
      20'h0714b: out <= 12'hb27;
      20'h0714c: out <= 12'hb27;
      20'h0714d: out <= 12'hb27;
      20'h0714e: out <= 12'hb27;
      20'h0714f: out <= 12'hb27;
      20'h07150: out <= 12'hb27;
      20'h07151: out <= 12'hb27;
      20'h07152: out <= 12'hb27;
      20'h07153: out <= 12'hb27;
      20'h07154: out <= 12'h603;
      20'h07155: out <= 12'h603;
      20'h07156: out <= 12'h603;
      20'h07157: out <= 12'h603;
      20'h07158: out <= 12'h603;
      20'h07159: out <= 12'h603;
      20'h0715a: out <= 12'h603;
      20'h0715b: out <= 12'h603;
      20'h0715c: out <= 12'h603;
      20'h0715d: out <= 12'h603;
      20'h0715e: out <= 12'h603;
      20'h0715f: out <= 12'h603;
      20'h07160: out <= 12'h603;
      20'h07161: out <= 12'h603;
      20'h07162: out <= 12'h603;
      20'h07163: out <= 12'h603;
      20'h07164: out <= 12'h603;
      20'h07165: out <= 12'h603;
      20'h07166: out <= 12'h603;
      20'h07167: out <= 12'h603;
      20'h07168: out <= 12'h603;
      20'h07169: out <= 12'h603;
      20'h0716a: out <= 12'h603;
      20'h0716b: out <= 12'h603;
      20'h0716c: out <= 12'h603;
      20'h0716d: out <= 12'h603;
      20'h0716e: out <= 12'h603;
      20'h0716f: out <= 12'h603;
      20'h07170: out <= 12'h603;
      20'h07171: out <= 12'h603;
      20'h07172: out <= 12'h603;
      20'h07173: out <= 12'h603;
      20'h07174: out <= 12'h603;
      20'h07175: out <= 12'h603;
      20'h07176: out <= 12'h603;
      20'h07177: out <= 12'h603;
      20'h07178: out <= 12'h603;
      20'h07179: out <= 12'h603;
      20'h0717a: out <= 12'h603;
      20'h0717b: out <= 12'h603;
      20'h0717c: out <= 12'h603;
      20'h0717d: out <= 12'h603;
      20'h0717e: out <= 12'h603;
      20'h0717f: out <= 12'h603;
      20'h07180: out <= 12'hb27;
      20'h07181: out <= 12'hb27;
      20'h07182: out <= 12'hb27;
      20'h07183: out <= 12'hb27;
      20'h07184: out <= 12'hb27;
      20'h07185: out <= 12'hb27;
      20'h07186: out <= 12'hb27;
      20'h07187: out <= 12'hb27;
      20'h07188: out <= 12'h000;
      20'h07189: out <= 12'h000;
      20'h0718a: out <= 12'h000;
      20'h0718b: out <= 12'h000;
      20'h0718c: out <= 12'h000;
      20'h0718d: out <= 12'h000;
      20'h0718e: out <= 12'h000;
      20'h0718f: out <= 12'h000;
      20'h07190: out <= 12'h777;
      20'h07191: out <= 12'h555;
      20'h07192: out <= 12'h555;
      20'h07193: out <= 12'h555;
      20'h07194: out <= 12'h555;
      20'h07195: out <= 12'h555;
      20'h07196: out <= 12'h555;
      20'h07197: out <= 12'h555;
      20'h07198: out <= 12'h555;
      20'h07199: out <= 12'h555;
      20'h0719a: out <= 12'h555;
      20'h0719b: out <= 12'h555;
      20'h0719c: out <= 12'h555;
      20'h0719d: out <= 12'h555;
      20'h0719e: out <= 12'h555;
      20'h0719f: out <= 12'h777;
      20'h071a0: out <= 12'h000;
      20'h071a1: out <= 12'h000;
      20'h071a2: out <= 12'h000;
      20'h071a3: out <= 12'h000;
      20'h071a4: out <= 12'h000;
      20'h071a5: out <= 12'h000;
      20'h071a6: out <= 12'h000;
      20'h071a7: out <= 12'h000;
      20'h071a8: out <= 12'h000;
      20'h071a9: out <= 12'h000;
      20'h071aa: out <= 12'h000;
      20'h071ab: out <= 12'h000;
      20'h071ac: out <= 12'h000;
      20'h071ad: out <= 12'h000;
      20'h071ae: out <= 12'h000;
      20'h071af: out <= 12'h000;
      20'h071b0: out <= 12'h000;
      20'h071b1: out <= 12'h000;
      20'h071b2: out <= 12'h000;
      20'h071b3: out <= 12'h000;
      20'h071b4: out <= 12'h000;
      20'h071b5: out <= 12'h000;
      20'h071b6: out <= 12'h000;
      20'h071b7: out <= 12'h000;
      20'h071b8: out <= 12'h000;
      20'h071b9: out <= 12'h000;
      20'h071ba: out <= 12'h000;
      20'h071bb: out <= 12'h000;
      20'h071bc: out <= 12'h000;
      20'h071bd: out <= 12'h000;
      20'h071be: out <= 12'h000;
      20'h071bf: out <= 12'h000;
      20'h071c0: out <= 12'h222;
      20'h071c1: out <= 12'h666;
      20'h071c2: out <= 12'hbbb;
      20'h071c3: out <= 12'hbbb;
      20'h071c4: out <= 12'h666;
      20'h071c5: out <= 12'h666;
      20'h071c6: out <= 12'hbbb;
      20'h071c7: out <= 12'hbbb;
      20'h071c8: out <= 12'h666;
      20'h071c9: out <= 12'hbbb;
      20'h071ca: out <= 12'hbbb;
      20'h071cb: out <= 12'hbbb;
      20'h071cc: out <= 12'hbbb;
      20'h071cd: out <= 12'hbbb;
      20'h071ce: out <= 12'hbbb;
      20'h071cf: out <= 12'hbbb;
      20'h071d0: out <= 12'h000;
      20'h071d1: out <= 12'h666;
      20'h071d2: out <= 12'hbbb;
      20'h071d3: out <= 12'hbbb;
      20'h071d4: out <= 12'h666;
      20'h071d5: out <= 12'h666;
      20'h071d6: out <= 12'hbbb;
      20'h071d7: out <= 12'hbbb;
      20'h071d8: out <= 12'h666;
      20'h071d9: out <= 12'hbbb;
      20'h071da: out <= 12'hbbb;
      20'h071db: out <= 12'hbbb;
      20'h071dc: out <= 12'hbbb;
      20'h071dd: out <= 12'hbbb;
      20'h071de: out <= 12'hbbb;
      20'h071df: out <= 12'hbbb;
      20'h071e0: out <= 12'h222;
      20'h071e1: out <= 12'h222;
      20'h071e2: out <= 12'h666;
      20'h071e3: out <= 12'h666;
      20'h071e4: out <= 12'h666;
      20'h071e5: out <= 12'hfff;
      20'h071e6: out <= 12'h666;
      20'h071e7: out <= 12'hfff;
      20'h071e8: out <= 12'hfff;
      20'h071e9: out <= 12'hbbb;
      20'h071ea: out <= 12'h666;
      20'h071eb: out <= 12'h666;
      20'h071ec: out <= 12'h666;
      20'h071ed: out <= 12'h666;
      20'h071ee: out <= 12'h666;
      20'h071ef: out <= 12'h222;
      20'h071f0: out <= 12'h000;
      20'h071f1: out <= 12'h000;
      20'h071f2: out <= 12'h666;
      20'h071f3: out <= 12'hbbb;
      20'h071f4: out <= 12'h666;
      20'h071f5: out <= 12'hfff;
      20'h071f6: out <= 12'h666;
      20'h071f7: out <= 12'hfff;
      20'h071f8: out <= 12'hfff;
      20'h071f9: out <= 12'hbbb;
      20'h071fa: out <= 12'h666;
      20'h071fb: out <= 12'h666;
      20'h071fc: out <= 12'h666;
      20'h071fd: out <= 12'hbbb;
      20'h071fe: out <= 12'h666;
      20'h071ff: out <= 12'h000;
      20'h07200: out <= 12'hbbb;
      20'h07201: out <= 12'hbbb;
      20'h07202: out <= 12'hbbb;
      20'h07203: out <= 12'hbbb;
      20'h07204: out <= 12'hbbb;
      20'h07205: out <= 12'hbbb;
      20'h07206: out <= 12'hbbb;
      20'h07207: out <= 12'h666;
      20'h07208: out <= 12'hbbb;
      20'h07209: out <= 12'hbbb;
      20'h0720a: out <= 12'h666;
      20'h0720b: out <= 12'h666;
      20'h0720c: out <= 12'hbbb;
      20'h0720d: out <= 12'hbbb;
      20'h0720e: out <= 12'h666;
      20'h0720f: out <= 12'h222;
      20'h07210: out <= 12'hbbb;
      20'h07211: out <= 12'hbbb;
      20'h07212: out <= 12'hbbb;
      20'h07213: out <= 12'hbbb;
      20'h07214: out <= 12'hbbb;
      20'h07215: out <= 12'hbbb;
      20'h07216: out <= 12'hbbb;
      20'h07217: out <= 12'h666;
      20'h07218: out <= 12'hbbb;
      20'h07219: out <= 12'hbbb;
      20'h0721a: out <= 12'h666;
      20'h0721b: out <= 12'h666;
      20'h0721c: out <= 12'hbbb;
      20'h0721d: out <= 12'hbbb;
      20'h0721e: out <= 12'h666;
      20'h0721f: out <= 12'h000;
      20'h07220: out <= 12'h222;
      20'h07221: out <= 12'h222;
      20'h07222: out <= 12'h222;
      20'h07223: out <= 12'hbbb;
      20'h07224: out <= 12'h666;
      20'h07225: out <= 12'hfff;
      20'h07226: out <= 12'hbbb;
      20'h07227: out <= 12'h666;
      20'h07228: out <= 12'h666;
      20'h07229: out <= 12'h666;
      20'h0722a: out <= 12'h666;
      20'h0722b: out <= 12'h666;
      20'h0722c: out <= 12'h666;
      20'h0722d: out <= 12'hbbb;
      20'h0722e: out <= 12'h222;
      20'h0722f: out <= 12'h222;
      20'h07230: out <= 12'h000;
      20'h07231: out <= 12'h000;
      20'h07232: out <= 12'h000;
      20'h07233: out <= 12'h666;
      20'h07234: out <= 12'h666;
      20'h07235: out <= 12'hfff;
      20'h07236: out <= 12'hbbb;
      20'h07237: out <= 12'h666;
      20'h07238: out <= 12'h666;
      20'h07239: out <= 12'h666;
      20'h0723a: out <= 12'h666;
      20'h0723b: out <= 12'h666;
      20'h0723c: out <= 12'h666;
      20'h0723d: out <= 12'h666;
      20'h0723e: out <= 12'h000;
      20'h0723f: out <= 12'h000;
      20'h07240: out <= 12'h603;
      20'h07241: out <= 12'h603;
      20'h07242: out <= 12'h603;
      20'h07243: out <= 12'h603;
      20'h07244: out <= 12'h603;
      20'h07245: out <= 12'h603;
      20'h07246: out <= 12'h603;
      20'h07247: out <= 12'h603;
      20'h07248: out <= 12'h603;
      20'h07249: out <= 12'h603;
      20'h0724a: out <= 12'h603;
      20'h0724b: out <= 12'h603;
      20'h0724c: out <= 12'hee9;
      20'h0724d: out <= 12'hee9;
      20'h0724e: out <= 12'hee9;
      20'h0724f: out <= 12'hee9;
      20'h07250: out <= 12'hee9;
      20'h07251: out <= 12'hee9;
      20'h07252: out <= 12'hee9;
      20'h07253: out <= 12'hb27;
      20'h07254: out <= 12'h603;
      20'h07255: out <= 12'h603;
      20'h07256: out <= 12'h603;
      20'h07257: out <= 12'h603;
      20'h07258: out <= 12'h603;
      20'h07259: out <= 12'h603;
      20'h0725a: out <= 12'h603;
      20'h0725b: out <= 12'h603;
      20'h0725c: out <= 12'h603;
      20'h0725d: out <= 12'h603;
      20'h0725e: out <= 12'h603;
      20'h0725f: out <= 12'h603;
      20'h07260: out <= 12'h603;
      20'h07261: out <= 12'h603;
      20'h07262: out <= 12'h603;
      20'h07263: out <= 12'h603;
      20'h07264: out <= 12'hee9;
      20'h07265: out <= 12'hee9;
      20'h07266: out <= 12'hee9;
      20'h07267: out <= 12'hee9;
      20'h07268: out <= 12'hee9;
      20'h07269: out <= 12'hee9;
      20'h0726a: out <= 12'hee9;
      20'h0726b: out <= 12'hb27;
      20'h0726c: out <= 12'h603;
      20'h0726d: out <= 12'h603;
      20'h0726e: out <= 12'h603;
      20'h0726f: out <= 12'h603;
      20'h07270: out <= 12'h603;
      20'h07271: out <= 12'h603;
      20'h07272: out <= 12'h603;
      20'h07273: out <= 12'h603;
      20'h07274: out <= 12'h603;
      20'h07275: out <= 12'h603;
      20'h07276: out <= 12'h603;
      20'h07277: out <= 12'h603;
      20'h07278: out <= 12'h603;
      20'h07279: out <= 12'h603;
      20'h0727a: out <= 12'h603;
      20'h0727b: out <= 12'h603;
      20'h0727c: out <= 12'h603;
      20'h0727d: out <= 12'h603;
      20'h0727e: out <= 12'h603;
      20'h0727f: out <= 12'h603;
      20'h07280: out <= 12'h603;
      20'h07281: out <= 12'h603;
      20'h07282: out <= 12'h603;
      20'h07283: out <= 12'h603;
      20'h07284: out <= 12'h603;
      20'h07285: out <= 12'h603;
      20'h07286: out <= 12'h603;
      20'h07287: out <= 12'h603;
      20'h07288: out <= 12'h603;
      20'h07289: out <= 12'h603;
      20'h0728a: out <= 12'h603;
      20'h0728b: out <= 12'h603;
      20'h0728c: out <= 12'h603;
      20'h0728d: out <= 12'h603;
      20'h0728e: out <= 12'h603;
      20'h0728f: out <= 12'h603;
      20'h07290: out <= 12'h603;
      20'h07291: out <= 12'h603;
      20'h07292: out <= 12'h603;
      20'h07293: out <= 12'h603;
      20'h07294: out <= 12'h603;
      20'h07295: out <= 12'h603;
      20'h07296: out <= 12'h603;
      20'h07297: out <= 12'h603;
      20'h07298: out <= 12'hee9;
      20'h07299: out <= 12'hee9;
      20'h0729a: out <= 12'hee9;
      20'h0729b: out <= 12'hee9;
      20'h0729c: out <= 12'hee9;
      20'h0729d: out <= 12'hee9;
      20'h0729e: out <= 12'hee9;
      20'h0729f: out <= 12'hb27;
      20'h072a0: out <= 12'h000;
      20'h072a1: out <= 12'h000;
      20'h072a2: out <= 12'h000;
      20'h072a3: out <= 12'h000;
      20'h072a4: out <= 12'h000;
      20'h072a5: out <= 12'h000;
      20'h072a6: out <= 12'h000;
      20'h072a7: out <= 12'h000;
      20'h072a8: out <= 12'h777;
      20'h072a9: out <= 12'h555;
      20'h072aa: out <= 12'h555;
      20'h072ab: out <= 12'h555;
      20'h072ac: out <= 12'h555;
      20'h072ad: out <= 12'h555;
      20'h072ae: out <= 12'h555;
      20'h072af: out <= 12'h555;
      20'h072b0: out <= 12'h555;
      20'h072b1: out <= 12'h555;
      20'h072b2: out <= 12'h555;
      20'h072b3: out <= 12'h555;
      20'h072b4: out <= 12'h555;
      20'h072b5: out <= 12'h555;
      20'h072b6: out <= 12'h555;
      20'h072b7: out <= 12'h777;
      20'h072b8: out <= 12'h000;
      20'h072b9: out <= 12'h000;
      20'h072ba: out <= 12'h000;
      20'h072bb: out <= 12'h000;
      20'h072bc: out <= 12'h000;
      20'h072bd: out <= 12'h000;
      20'h072be: out <= 12'h000;
      20'h072bf: out <= 12'h000;
      20'h072c0: out <= 12'hfa9;
      20'h072c1: out <= 12'hfa9;
      20'h072c2: out <= 12'hfa9;
      20'h072c3: out <= 12'hfa9;
      20'h072c4: out <= 12'hfa9;
      20'h072c5: out <= 12'hfa9;
      20'h072c6: out <= 12'hfa9;
      20'h072c7: out <= 12'hfa9;
      20'h072c8: out <= 12'hf76;
      20'h072c9: out <= 12'hf76;
      20'h072ca: out <= 12'hf76;
      20'h072cb: out <= 12'hf76;
      20'h072cc: out <= 12'hf76;
      20'h072cd: out <= 12'hf76;
      20'h072ce: out <= 12'hf76;
      20'h072cf: out <= 12'hf76;
      20'h072d0: out <= 12'h000;
      20'h072d1: out <= 12'h000;
      20'h072d2: out <= 12'h000;
      20'h072d3: out <= 12'h000;
      20'h072d4: out <= 12'h000;
      20'h072d5: out <= 12'h000;
      20'h072d6: out <= 12'h000;
      20'h072d7: out <= 12'h000;
      20'h072d8: out <= 12'h222;
      20'h072d9: out <= 12'h666;
      20'h072da: out <= 12'h666;
      20'h072db: out <= 12'h666;
      20'h072dc: out <= 12'h666;
      20'h072dd: out <= 12'h666;
      20'h072de: out <= 12'h666;
      20'h072df: out <= 12'h666;
      20'h072e0: out <= 12'h666;
      20'h072e1: out <= 12'h666;
      20'h072e2: out <= 12'h666;
      20'h072e3: out <= 12'h666;
      20'h072e4: out <= 12'h666;
      20'h072e5: out <= 12'h666;
      20'h072e6: out <= 12'h666;
      20'h072e7: out <= 12'h666;
      20'h072e8: out <= 12'h000;
      20'h072e9: out <= 12'h666;
      20'h072ea: out <= 12'h666;
      20'h072eb: out <= 12'h666;
      20'h072ec: out <= 12'h666;
      20'h072ed: out <= 12'h666;
      20'h072ee: out <= 12'h666;
      20'h072ef: out <= 12'h666;
      20'h072f0: out <= 12'h666;
      20'h072f1: out <= 12'h666;
      20'h072f2: out <= 12'h666;
      20'h072f3: out <= 12'h666;
      20'h072f4: out <= 12'h666;
      20'h072f5: out <= 12'h666;
      20'h072f6: out <= 12'h666;
      20'h072f7: out <= 12'h666;
      20'h072f8: out <= 12'h222;
      20'h072f9: out <= 12'h222;
      20'h072fa: out <= 12'h222;
      20'h072fb: out <= 12'hbbb;
      20'h072fc: out <= 12'h666;
      20'h072fd: out <= 12'hfff;
      20'h072fe: out <= 12'h666;
      20'h072ff: out <= 12'hfff;
      20'h07300: out <= 12'hbbb;
      20'h07301: out <= 12'hbbb;
      20'h07302: out <= 12'h666;
      20'h07303: out <= 12'h666;
      20'h07304: out <= 12'h666;
      20'h07305: out <= 12'hbbb;
      20'h07306: out <= 12'h222;
      20'h07307: out <= 12'h222;
      20'h07308: out <= 12'h000;
      20'h07309: out <= 12'h000;
      20'h0730a: out <= 12'h000;
      20'h0730b: out <= 12'h666;
      20'h0730c: out <= 12'h666;
      20'h0730d: out <= 12'hfff;
      20'h0730e: out <= 12'h666;
      20'h0730f: out <= 12'hfff;
      20'h07310: out <= 12'hbbb;
      20'h07311: out <= 12'hbbb;
      20'h07312: out <= 12'h666;
      20'h07313: out <= 12'h666;
      20'h07314: out <= 12'h666;
      20'h07315: out <= 12'h666;
      20'h07316: out <= 12'h000;
      20'h07317: out <= 12'h000;
      20'h07318: out <= 12'h666;
      20'h07319: out <= 12'h666;
      20'h0731a: out <= 12'h666;
      20'h0731b: out <= 12'h666;
      20'h0731c: out <= 12'h666;
      20'h0731d: out <= 12'h666;
      20'h0731e: out <= 12'h666;
      20'h0731f: out <= 12'h666;
      20'h07320: out <= 12'h666;
      20'h07321: out <= 12'h666;
      20'h07322: out <= 12'h666;
      20'h07323: out <= 12'h666;
      20'h07324: out <= 12'h666;
      20'h07325: out <= 12'h666;
      20'h07326: out <= 12'h666;
      20'h07327: out <= 12'h222;
      20'h07328: out <= 12'h666;
      20'h07329: out <= 12'h666;
      20'h0732a: out <= 12'h666;
      20'h0732b: out <= 12'h666;
      20'h0732c: out <= 12'h666;
      20'h0732d: out <= 12'h666;
      20'h0732e: out <= 12'h666;
      20'h0732f: out <= 12'h666;
      20'h07330: out <= 12'h666;
      20'h07331: out <= 12'h666;
      20'h07332: out <= 12'h666;
      20'h07333: out <= 12'h666;
      20'h07334: out <= 12'h666;
      20'h07335: out <= 12'h666;
      20'h07336: out <= 12'h666;
      20'h07337: out <= 12'h000;
      20'h07338: out <= 12'h222;
      20'h07339: out <= 12'h222;
      20'h0733a: out <= 12'h666;
      20'h0733b: out <= 12'h666;
      20'h0733c: out <= 12'h666;
      20'h0733d: out <= 12'hfff;
      20'h0733e: out <= 12'h666;
      20'h0733f: out <= 12'hbbb;
      20'h07340: out <= 12'hfff;
      20'h07341: out <= 12'hbbb;
      20'h07342: out <= 12'h666;
      20'h07343: out <= 12'h666;
      20'h07344: out <= 12'h666;
      20'h07345: out <= 12'h666;
      20'h07346: out <= 12'h666;
      20'h07347: out <= 12'h222;
      20'h07348: out <= 12'h000;
      20'h07349: out <= 12'h000;
      20'h0734a: out <= 12'h666;
      20'h0734b: out <= 12'hbbb;
      20'h0734c: out <= 12'h666;
      20'h0734d: out <= 12'hfff;
      20'h0734e: out <= 12'h666;
      20'h0734f: out <= 12'hbbb;
      20'h07350: out <= 12'hfff;
      20'h07351: out <= 12'hbbb;
      20'h07352: out <= 12'h666;
      20'h07353: out <= 12'h666;
      20'h07354: out <= 12'h666;
      20'h07355: out <= 12'hbbb;
      20'h07356: out <= 12'h666;
      20'h07357: out <= 12'h000;
      20'h07358: out <= 12'h603;
      20'h07359: out <= 12'h603;
      20'h0735a: out <= 12'h603;
      20'h0735b: out <= 12'h603;
      20'h0735c: out <= 12'h603;
      20'h0735d: out <= 12'h603;
      20'h0735e: out <= 12'h603;
      20'h0735f: out <= 12'h603;
      20'h07360: out <= 12'h603;
      20'h07361: out <= 12'h603;
      20'h07362: out <= 12'h603;
      20'h07363: out <= 12'h603;
      20'h07364: out <= 12'hee9;
      20'h07365: out <= 12'hf87;
      20'h07366: out <= 12'hf87;
      20'h07367: out <= 12'hf87;
      20'h07368: out <= 12'hf87;
      20'h07369: out <= 12'hf87;
      20'h0736a: out <= 12'hf87;
      20'h0736b: out <= 12'hb27;
      20'h0736c: out <= 12'h603;
      20'h0736d: out <= 12'h603;
      20'h0736e: out <= 12'h603;
      20'h0736f: out <= 12'h603;
      20'h07370: out <= 12'h603;
      20'h07371: out <= 12'h603;
      20'h07372: out <= 12'h603;
      20'h07373: out <= 12'h603;
      20'h07374: out <= 12'h603;
      20'h07375: out <= 12'h603;
      20'h07376: out <= 12'h603;
      20'h07377: out <= 12'h603;
      20'h07378: out <= 12'h603;
      20'h07379: out <= 12'h603;
      20'h0737a: out <= 12'h603;
      20'h0737b: out <= 12'h603;
      20'h0737c: out <= 12'hee9;
      20'h0737d: out <= 12'hf87;
      20'h0737e: out <= 12'hf87;
      20'h0737f: out <= 12'hf87;
      20'h07380: out <= 12'hf87;
      20'h07381: out <= 12'hf87;
      20'h07382: out <= 12'hf87;
      20'h07383: out <= 12'hb27;
      20'h07384: out <= 12'h603;
      20'h07385: out <= 12'h603;
      20'h07386: out <= 12'h603;
      20'h07387: out <= 12'h603;
      20'h07388: out <= 12'h603;
      20'h07389: out <= 12'h603;
      20'h0738a: out <= 12'h603;
      20'h0738b: out <= 12'h603;
      20'h0738c: out <= 12'h603;
      20'h0738d: out <= 12'h603;
      20'h0738e: out <= 12'h603;
      20'h0738f: out <= 12'h603;
      20'h07390: out <= 12'h603;
      20'h07391: out <= 12'h603;
      20'h07392: out <= 12'h603;
      20'h07393: out <= 12'h603;
      20'h07394: out <= 12'h603;
      20'h07395: out <= 12'h603;
      20'h07396: out <= 12'h603;
      20'h07397: out <= 12'h603;
      20'h07398: out <= 12'h603;
      20'h07399: out <= 12'h603;
      20'h0739a: out <= 12'h603;
      20'h0739b: out <= 12'h603;
      20'h0739c: out <= 12'h603;
      20'h0739d: out <= 12'h603;
      20'h0739e: out <= 12'h603;
      20'h0739f: out <= 12'h603;
      20'h073a0: out <= 12'h603;
      20'h073a1: out <= 12'h603;
      20'h073a2: out <= 12'h603;
      20'h073a3: out <= 12'h603;
      20'h073a4: out <= 12'h603;
      20'h073a5: out <= 12'h603;
      20'h073a6: out <= 12'h603;
      20'h073a7: out <= 12'h603;
      20'h073a8: out <= 12'h603;
      20'h073a9: out <= 12'h603;
      20'h073aa: out <= 12'h603;
      20'h073ab: out <= 12'h603;
      20'h073ac: out <= 12'h603;
      20'h073ad: out <= 12'h603;
      20'h073ae: out <= 12'h603;
      20'h073af: out <= 12'h603;
      20'h073b0: out <= 12'hee9;
      20'h073b1: out <= 12'hf87;
      20'h073b2: out <= 12'hf87;
      20'h073b3: out <= 12'hf87;
      20'h073b4: out <= 12'hf87;
      20'h073b5: out <= 12'hf87;
      20'h073b6: out <= 12'hf87;
      20'h073b7: out <= 12'hb27;
      20'h073b8: out <= 12'h000;
      20'h073b9: out <= 12'h000;
      20'h073ba: out <= 12'h000;
      20'h073bb: out <= 12'h000;
      20'h073bc: out <= 12'h000;
      20'h073bd: out <= 12'h000;
      20'h073be: out <= 12'h000;
      20'h073bf: out <= 12'h000;
      20'h073c0: out <= 12'h777;
      20'h073c1: out <= 12'h555;
      20'h073c2: out <= 12'h555;
      20'h073c3: out <= 12'h555;
      20'h073c4: out <= 12'h555;
      20'h073c5: out <= 12'h555;
      20'h073c6: out <= 12'h555;
      20'h073c7: out <= 12'h555;
      20'h073c8: out <= 12'h555;
      20'h073c9: out <= 12'h555;
      20'h073ca: out <= 12'h555;
      20'h073cb: out <= 12'h555;
      20'h073cc: out <= 12'h555;
      20'h073cd: out <= 12'h555;
      20'h073ce: out <= 12'h555;
      20'h073cf: out <= 12'h777;
      20'h073d0: out <= 12'h000;
      20'h073d1: out <= 12'h000;
      20'h073d2: out <= 12'hf87;
      20'h073d3: out <= 12'h000;
      20'h073d4: out <= 12'h000;
      20'h073d5: out <= 12'h000;
      20'h073d6: out <= 12'hf87;
      20'h073d7: out <= 12'h000;
      20'h073d8: out <= 12'hfa9;
      20'h073d9: out <= 12'hfa9;
      20'h073da: out <= 12'hfa9;
      20'h073db: out <= 12'hfa9;
      20'h073dc: out <= 12'hfa9;
      20'h073dd: out <= 12'hfa9;
      20'h073de: out <= 12'hfa9;
      20'h073df: out <= 12'hfa9;
      20'h073e0: out <= 12'hf76;
      20'h073e1: out <= 12'hf76;
      20'h073e2: out <= 12'hf76;
      20'h073e3: out <= 12'hf76;
      20'h073e4: out <= 12'hf76;
      20'h073e5: out <= 12'hf76;
      20'h073e6: out <= 12'hf76;
      20'h073e7: out <= 12'hf76;
      20'h073e8: out <= 12'h000;
      20'h073e9: out <= 12'h000;
      20'h073ea: out <= 12'h000;
      20'h073eb: out <= 12'h000;
      20'h073ec: out <= 12'h000;
      20'h073ed: out <= 12'h000;
      20'h073ee: out <= 12'h000;
      20'h073ef: out <= 12'h000;
      20'h073f0: out <= 12'h222;
      20'h073f1: out <= 12'h222;
      20'h073f2: out <= 12'h666;
      20'h073f3: out <= 12'h666;
      20'h073f4: out <= 12'h666;
      20'h073f5: out <= 12'h666;
      20'h073f6: out <= 12'h666;
      20'h073f7: out <= 12'h666;
      20'h073f8: out <= 12'h666;
      20'h073f9: out <= 12'h666;
      20'h073fa: out <= 12'h666;
      20'h073fb: out <= 12'h666;
      20'h073fc: out <= 12'h666;
      20'h073fd: out <= 12'h222;
      20'h073fe: out <= 12'h222;
      20'h073ff: out <= 12'h222;
      20'h07400: out <= 12'h000;
      20'h07401: out <= 12'h000;
      20'h07402: out <= 12'h666;
      20'h07403: out <= 12'h666;
      20'h07404: out <= 12'h666;
      20'h07405: out <= 12'h666;
      20'h07406: out <= 12'h666;
      20'h07407: out <= 12'h666;
      20'h07408: out <= 12'h666;
      20'h07409: out <= 12'h666;
      20'h0740a: out <= 12'h666;
      20'h0740b: out <= 12'h666;
      20'h0740c: out <= 12'h666;
      20'h0740d: out <= 12'h000;
      20'h0740e: out <= 12'h000;
      20'h0740f: out <= 12'h000;
      20'h07410: out <= 12'h222;
      20'h07411: out <= 12'h222;
      20'h07412: out <= 12'h666;
      20'h07413: out <= 12'h666;
      20'h07414: out <= 12'h666;
      20'h07415: out <= 12'hfff;
      20'h07416: out <= 12'h666;
      20'h07417: out <= 12'hbbb;
      20'h07418: out <= 12'hbbb;
      20'h07419: out <= 12'h666;
      20'h0741a: out <= 12'h666;
      20'h0741b: out <= 12'h666;
      20'h0741c: out <= 12'h666;
      20'h0741d: out <= 12'h666;
      20'h0741e: out <= 12'h666;
      20'h0741f: out <= 12'h222;
      20'h07420: out <= 12'h000;
      20'h07421: out <= 12'h000;
      20'h07422: out <= 12'h666;
      20'h07423: out <= 12'hbbb;
      20'h07424: out <= 12'h666;
      20'h07425: out <= 12'hfff;
      20'h07426: out <= 12'h666;
      20'h07427: out <= 12'hbbb;
      20'h07428: out <= 12'hbbb;
      20'h07429: out <= 12'h666;
      20'h0742a: out <= 12'h666;
      20'h0742b: out <= 12'h666;
      20'h0742c: out <= 12'h666;
      20'h0742d: out <= 12'hbbb;
      20'h0742e: out <= 12'h666;
      20'h0742f: out <= 12'h000;
      20'h07430: out <= 12'h222;
      20'h07431: out <= 12'h222;
      20'h07432: out <= 12'h222;
      20'h07433: out <= 12'h666;
      20'h07434: out <= 12'h666;
      20'h07435: out <= 12'h666;
      20'h07436: out <= 12'h666;
      20'h07437: out <= 12'h666;
      20'h07438: out <= 12'h666;
      20'h07439: out <= 12'h666;
      20'h0743a: out <= 12'h666;
      20'h0743b: out <= 12'h666;
      20'h0743c: out <= 12'h666;
      20'h0743d: out <= 12'h666;
      20'h0743e: out <= 12'h222;
      20'h0743f: out <= 12'h222;
      20'h07440: out <= 12'h000;
      20'h07441: out <= 12'h000;
      20'h07442: out <= 12'h000;
      20'h07443: out <= 12'h666;
      20'h07444: out <= 12'h666;
      20'h07445: out <= 12'h666;
      20'h07446: out <= 12'h666;
      20'h07447: out <= 12'h666;
      20'h07448: out <= 12'h666;
      20'h07449: out <= 12'h666;
      20'h0744a: out <= 12'h666;
      20'h0744b: out <= 12'h666;
      20'h0744c: out <= 12'h666;
      20'h0744d: out <= 12'h666;
      20'h0744e: out <= 12'h000;
      20'h0744f: out <= 12'h000;
      20'h07450: out <= 12'h222;
      20'h07451: out <= 12'h222;
      20'h07452: out <= 12'h222;
      20'h07453: out <= 12'hbbb;
      20'h07454: out <= 12'h666;
      20'h07455: out <= 12'hfff;
      20'h07456: out <= 12'h666;
      20'h07457: out <= 12'hbbb;
      20'h07458: out <= 12'hfff;
      20'h07459: out <= 12'hbbb;
      20'h0745a: out <= 12'h666;
      20'h0745b: out <= 12'h666;
      20'h0745c: out <= 12'h666;
      20'h0745d: out <= 12'hbbb;
      20'h0745e: out <= 12'h222;
      20'h0745f: out <= 12'h222;
      20'h07460: out <= 12'h000;
      20'h07461: out <= 12'h000;
      20'h07462: out <= 12'h000;
      20'h07463: out <= 12'h666;
      20'h07464: out <= 12'h666;
      20'h07465: out <= 12'hfff;
      20'h07466: out <= 12'h666;
      20'h07467: out <= 12'hbbb;
      20'h07468: out <= 12'hfff;
      20'h07469: out <= 12'hbbb;
      20'h0746a: out <= 12'h666;
      20'h0746b: out <= 12'h666;
      20'h0746c: out <= 12'h666;
      20'h0746d: out <= 12'h666;
      20'h0746e: out <= 12'h000;
      20'h0746f: out <= 12'h000;
      20'h07470: out <= 12'h603;
      20'h07471: out <= 12'h603;
      20'h07472: out <= 12'h603;
      20'h07473: out <= 12'h603;
      20'h07474: out <= 12'h603;
      20'h07475: out <= 12'h603;
      20'h07476: out <= 12'h603;
      20'h07477: out <= 12'h603;
      20'h07478: out <= 12'h603;
      20'h07479: out <= 12'h603;
      20'h0747a: out <= 12'h603;
      20'h0747b: out <= 12'h603;
      20'h0747c: out <= 12'hee9;
      20'h0747d: out <= 12'hf87;
      20'h0747e: out <= 12'hee9;
      20'h0747f: out <= 12'hee9;
      20'h07480: out <= 12'hee9;
      20'h07481: out <= 12'hb27;
      20'h07482: out <= 12'hf87;
      20'h07483: out <= 12'hb27;
      20'h07484: out <= 12'h603;
      20'h07485: out <= 12'h603;
      20'h07486: out <= 12'h603;
      20'h07487: out <= 12'h603;
      20'h07488: out <= 12'h603;
      20'h07489: out <= 12'h603;
      20'h0748a: out <= 12'h603;
      20'h0748b: out <= 12'h603;
      20'h0748c: out <= 12'h603;
      20'h0748d: out <= 12'h603;
      20'h0748e: out <= 12'h603;
      20'h0748f: out <= 12'h603;
      20'h07490: out <= 12'h603;
      20'h07491: out <= 12'h603;
      20'h07492: out <= 12'h603;
      20'h07493: out <= 12'h603;
      20'h07494: out <= 12'hee9;
      20'h07495: out <= 12'hf87;
      20'h07496: out <= 12'hee9;
      20'h07497: out <= 12'hee9;
      20'h07498: out <= 12'hee9;
      20'h07499: out <= 12'hb27;
      20'h0749a: out <= 12'hf87;
      20'h0749b: out <= 12'hb27;
      20'h0749c: out <= 12'h603;
      20'h0749d: out <= 12'h603;
      20'h0749e: out <= 12'h603;
      20'h0749f: out <= 12'h603;
      20'h074a0: out <= 12'h603;
      20'h074a1: out <= 12'h603;
      20'h074a2: out <= 12'h603;
      20'h074a3: out <= 12'h603;
      20'h074a4: out <= 12'h603;
      20'h074a5: out <= 12'h603;
      20'h074a6: out <= 12'h603;
      20'h074a7: out <= 12'h603;
      20'h074a8: out <= 12'h603;
      20'h074a9: out <= 12'h603;
      20'h074aa: out <= 12'h603;
      20'h074ab: out <= 12'h603;
      20'h074ac: out <= 12'h603;
      20'h074ad: out <= 12'h603;
      20'h074ae: out <= 12'h603;
      20'h074af: out <= 12'h603;
      20'h074b0: out <= 12'h603;
      20'h074b1: out <= 12'h603;
      20'h074b2: out <= 12'h603;
      20'h074b3: out <= 12'h603;
      20'h074b4: out <= 12'h603;
      20'h074b5: out <= 12'h603;
      20'h074b6: out <= 12'h603;
      20'h074b7: out <= 12'h603;
      20'h074b8: out <= 12'h603;
      20'h074b9: out <= 12'h603;
      20'h074ba: out <= 12'h603;
      20'h074bb: out <= 12'h603;
      20'h074bc: out <= 12'h603;
      20'h074bd: out <= 12'h603;
      20'h074be: out <= 12'h603;
      20'h074bf: out <= 12'h603;
      20'h074c0: out <= 12'h603;
      20'h074c1: out <= 12'h603;
      20'h074c2: out <= 12'h603;
      20'h074c3: out <= 12'h603;
      20'h074c4: out <= 12'h603;
      20'h074c5: out <= 12'h603;
      20'h074c6: out <= 12'h603;
      20'h074c7: out <= 12'h603;
      20'h074c8: out <= 12'hee9;
      20'h074c9: out <= 12'hf87;
      20'h074ca: out <= 12'hee9;
      20'h074cb: out <= 12'hee9;
      20'h074cc: out <= 12'hee9;
      20'h074cd: out <= 12'hb27;
      20'h074ce: out <= 12'hf87;
      20'h074cf: out <= 12'hb27;
      20'h074d0: out <= 12'h000;
      20'h074d1: out <= 12'h000;
      20'h074d2: out <= 12'h000;
      20'h074d3: out <= 12'h000;
      20'h074d4: out <= 12'h000;
      20'h074d5: out <= 12'h000;
      20'h074d6: out <= 12'h000;
      20'h074d7: out <= 12'h000;
      20'h074d8: out <= 12'h777;
      20'h074d9: out <= 12'h555;
      20'h074da: out <= 12'h555;
      20'h074db: out <= 12'h555;
      20'h074dc: out <= 12'h555;
      20'h074dd: out <= 12'h555;
      20'h074de: out <= 12'h555;
      20'h074df: out <= 12'h555;
      20'h074e0: out <= 12'h555;
      20'h074e1: out <= 12'h555;
      20'h074e2: out <= 12'h555;
      20'h074e3: out <= 12'h555;
      20'h074e4: out <= 12'h555;
      20'h074e5: out <= 12'h555;
      20'h074e6: out <= 12'h555;
      20'h074e7: out <= 12'h777;
      20'h074e8: out <= 12'h000;
      20'h074e9: out <= 12'h000;
      20'h074ea: out <= 12'h000;
      20'h074eb: out <= 12'hf87;
      20'h074ec: out <= 12'h000;
      20'h074ed: out <= 12'hf87;
      20'h074ee: out <= 12'h000;
      20'h074ef: out <= 12'h000;
      20'h074f0: out <= 12'hfa9;
      20'h074f1: out <= 12'hfa9;
      20'h074f2: out <= 12'hfa9;
      20'h074f3: out <= 12'hfa9;
      20'h074f4: out <= 12'hfa9;
      20'h074f5: out <= 12'hfa9;
      20'h074f6: out <= 12'hfa9;
      20'h074f7: out <= 12'hfa9;
      20'h074f8: out <= 12'hf76;
      20'h074f9: out <= 12'hf76;
      20'h074fa: out <= 12'hf76;
      20'h074fb: out <= 12'hf76;
      20'h074fc: out <= 12'hf76;
      20'h074fd: out <= 12'hf76;
      20'h074fe: out <= 12'hf76;
      20'h074ff: out <= 12'hf76;
      20'h07500: out <= 12'h000;
      20'h07501: out <= 12'h000;
      20'h07502: out <= 12'h000;
      20'h07503: out <= 12'h000;
      20'h07504: out <= 12'h000;
      20'h07505: out <= 12'h000;
      20'h07506: out <= 12'h000;
      20'h07507: out <= 12'h000;
      20'h07508: out <= 12'h222;
      20'h07509: out <= 12'h222;
      20'h0750a: out <= 12'h222;
      20'h0750b: out <= 12'h666;
      20'h0750c: out <= 12'h666;
      20'h0750d: out <= 12'h666;
      20'h0750e: out <= 12'h666;
      20'h0750f: out <= 12'h666;
      20'h07510: out <= 12'h666;
      20'h07511: out <= 12'h666;
      20'h07512: out <= 12'h666;
      20'h07513: out <= 12'h666;
      20'h07514: out <= 12'h222;
      20'h07515: out <= 12'h222;
      20'h07516: out <= 12'h222;
      20'h07517: out <= 12'h222;
      20'h07518: out <= 12'h000;
      20'h07519: out <= 12'h000;
      20'h0751a: out <= 12'h000;
      20'h0751b: out <= 12'h666;
      20'h0751c: out <= 12'h666;
      20'h0751d: out <= 12'h666;
      20'h0751e: out <= 12'h666;
      20'h0751f: out <= 12'h666;
      20'h07520: out <= 12'h666;
      20'h07521: out <= 12'h666;
      20'h07522: out <= 12'h666;
      20'h07523: out <= 12'h666;
      20'h07524: out <= 12'h000;
      20'h07525: out <= 12'h000;
      20'h07526: out <= 12'h000;
      20'h07527: out <= 12'h000;
      20'h07528: out <= 12'h222;
      20'h07529: out <= 12'h222;
      20'h0752a: out <= 12'h222;
      20'h0752b: out <= 12'hbbb;
      20'h0752c: out <= 12'h666;
      20'h0752d: out <= 12'hfff;
      20'h0752e: out <= 12'hfff;
      20'h0752f: out <= 12'h666;
      20'h07530: out <= 12'h666;
      20'h07531: out <= 12'h666;
      20'h07532: out <= 12'h666;
      20'h07533: out <= 12'h666;
      20'h07534: out <= 12'h666;
      20'h07535: out <= 12'hbbb;
      20'h07536: out <= 12'h222;
      20'h07537: out <= 12'h222;
      20'h07538: out <= 12'h000;
      20'h07539: out <= 12'h000;
      20'h0753a: out <= 12'h000;
      20'h0753b: out <= 12'h666;
      20'h0753c: out <= 12'h666;
      20'h0753d: out <= 12'hfff;
      20'h0753e: out <= 12'hfff;
      20'h0753f: out <= 12'h666;
      20'h07540: out <= 12'h666;
      20'h07541: out <= 12'h666;
      20'h07542: out <= 12'h666;
      20'h07543: out <= 12'h666;
      20'h07544: out <= 12'h666;
      20'h07545: out <= 12'h666;
      20'h07546: out <= 12'h000;
      20'h07547: out <= 12'h000;
      20'h07548: out <= 12'h222;
      20'h07549: out <= 12'h222;
      20'h0754a: out <= 12'h222;
      20'h0754b: out <= 12'h222;
      20'h0754c: out <= 12'h666;
      20'h0754d: out <= 12'h666;
      20'h0754e: out <= 12'h666;
      20'h0754f: out <= 12'h666;
      20'h07550: out <= 12'h666;
      20'h07551: out <= 12'h666;
      20'h07552: out <= 12'h666;
      20'h07553: out <= 12'h666;
      20'h07554: out <= 12'h666;
      20'h07555: out <= 12'h222;
      20'h07556: out <= 12'h222;
      20'h07557: out <= 12'h222;
      20'h07558: out <= 12'h000;
      20'h07559: out <= 12'h000;
      20'h0755a: out <= 12'h000;
      20'h0755b: out <= 12'h000;
      20'h0755c: out <= 12'h666;
      20'h0755d: out <= 12'h666;
      20'h0755e: out <= 12'h666;
      20'h0755f: out <= 12'h666;
      20'h07560: out <= 12'h666;
      20'h07561: out <= 12'h666;
      20'h07562: out <= 12'h666;
      20'h07563: out <= 12'h666;
      20'h07564: out <= 12'h666;
      20'h07565: out <= 12'h000;
      20'h07566: out <= 12'h000;
      20'h07567: out <= 12'h000;
      20'h07568: out <= 12'h222;
      20'h07569: out <= 12'h222;
      20'h0756a: out <= 12'h666;
      20'h0756b: out <= 12'h666;
      20'h0756c: out <= 12'h666;
      20'h0756d: out <= 12'hfff;
      20'h0756e: out <= 12'h666;
      20'h0756f: out <= 12'hbbb;
      20'h07570: out <= 12'hfff;
      20'h07571: out <= 12'hbbb;
      20'h07572: out <= 12'h666;
      20'h07573: out <= 12'h666;
      20'h07574: out <= 12'h666;
      20'h07575: out <= 12'h666;
      20'h07576: out <= 12'h666;
      20'h07577: out <= 12'h222;
      20'h07578: out <= 12'h000;
      20'h07579: out <= 12'h000;
      20'h0757a: out <= 12'h666;
      20'h0757b: out <= 12'hbbb;
      20'h0757c: out <= 12'h666;
      20'h0757d: out <= 12'hfff;
      20'h0757e: out <= 12'h666;
      20'h0757f: out <= 12'hbbb;
      20'h07580: out <= 12'hfff;
      20'h07581: out <= 12'hbbb;
      20'h07582: out <= 12'h666;
      20'h07583: out <= 12'h666;
      20'h07584: out <= 12'h666;
      20'h07585: out <= 12'hbbb;
      20'h07586: out <= 12'h666;
      20'h07587: out <= 12'h000;
      20'h07588: out <= 12'h603;
      20'h07589: out <= 12'h603;
      20'h0758a: out <= 12'h603;
      20'h0758b: out <= 12'h603;
      20'h0758c: out <= 12'h603;
      20'h0758d: out <= 12'h603;
      20'h0758e: out <= 12'h603;
      20'h0758f: out <= 12'h603;
      20'h07590: out <= 12'h603;
      20'h07591: out <= 12'h603;
      20'h07592: out <= 12'h603;
      20'h07593: out <= 12'h603;
      20'h07594: out <= 12'hee9;
      20'h07595: out <= 12'hf87;
      20'h07596: out <= 12'hee9;
      20'h07597: out <= 12'hf87;
      20'h07598: out <= 12'hf87;
      20'h07599: out <= 12'hb27;
      20'h0759a: out <= 12'hf87;
      20'h0759b: out <= 12'hb27;
      20'h0759c: out <= 12'h603;
      20'h0759d: out <= 12'h603;
      20'h0759e: out <= 12'h603;
      20'h0759f: out <= 12'h603;
      20'h075a0: out <= 12'h603;
      20'h075a1: out <= 12'h603;
      20'h075a2: out <= 12'h603;
      20'h075a3: out <= 12'h603;
      20'h075a4: out <= 12'h603;
      20'h075a5: out <= 12'h603;
      20'h075a6: out <= 12'h603;
      20'h075a7: out <= 12'h603;
      20'h075a8: out <= 12'h603;
      20'h075a9: out <= 12'h603;
      20'h075aa: out <= 12'h603;
      20'h075ab: out <= 12'h603;
      20'h075ac: out <= 12'hee9;
      20'h075ad: out <= 12'hf87;
      20'h075ae: out <= 12'hee9;
      20'h075af: out <= 12'hf87;
      20'h075b0: out <= 12'hf87;
      20'h075b1: out <= 12'hb27;
      20'h075b2: out <= 12'hf87;
      20'h075b3: out <= 12'hb27;
      20'h075b4: out <= 12'h603;
      20'h075b5: out <= 12'h603;
      20'h075b6: out <= 12'h603;
      20'h075b7: out <= 12'h603;
      20'h075b8: out <= 12'h603;
      20'h075b9: out <= 12'h603;
      20'h075ba: out <= 12'h603;
      20'h075bb: out <= 12'h603;
      20'h075bc: out <= 12'h603;
      20'h075bd: out <= 12'h603;
      20'h075be: out <= 12'h603;
      20'h075bf: out <= 12'h603;
      20'h075c0: out <= 12'h603;
      20'h075c1: out <= 12'h603;
      20'h075c2: out <= 12'h603;
      20'h075c3: out <= 12'h603;
      20'h075c4: out <= 12'h603;
      20'h075c5: out <= 12'h603;
      20'h075c6: out <= 12'h603;
      20'h075c7: out <= 12'h603;
      20'h075c8: out <= 12'h603;
      20'h075c9: out <= 12'h603;
      20'h075ca: out <= 12'h603;
      20'h075cb: out <= 12'h603;
      20'h075cc: out <= 12'h603;
      20'h075cd: out <= 12'h603;
      20'h075ce: out <= 12'h603;
      20'h075cf: out <= 12'h603;
      20'h075d0: out <= 12'h603;
      20'h075d1: out <= 12'h603;
      20'h075d2: out <= 12'h603;
      20'h075d3: out <= 12'h603;
      20'h075d4: out <= 12'h603;
      20'h075d5: out <= 12'h603;
      20'h075d6: out <= 12'h603;
      20'h075d7: out <= 12'h603;
      20'h075d8: out <= 12'h603;
      20'h075d9: out <= 12'h603;
      20'h075da: out <= 12'h603;
      20'h075db: out <= 12'h603;
      20'h075dc: out <= 12'h603;
      20'h075dd: out <= 12'h603;
      20'h075de: out <= 12'h603;
      20'h075df: out <= 12'h603;
      20'h075e0: out <= 12'hee9;
      20'h075e1: out <= 12'hf87;
      20'h075e2: out <= 12'hee9;
      20'h075e3: out <= 12'hf87;
      20'h075e4: out <= 12'hf87;
      20'h075e5: out <= 12'hb27;
      20'h075e6: out <= 12'hf87;
      20'h075e7: out <= 12'hb27;
      20'h075e8: out <= 12'h000;
      20'h075e9: out <= 12'h000;
      20'h075ea: out <= 12'h000;
      20'h075eb: out <= 12'h000;
      20'h075ec: out <= 12'h000;
      20'h075ed: out <= 12'h000;
      20'h075ee: out <= 12'h000;
      20'h075ef: out <= 12'h000;
      20'h075f0: out <= 12'h777;
      20'h075f1: out <= 12'h555;
      20'h075f2: out <= 12'h555;
      20'h075f3: out <= 12'h555;
      20'h075f4: out <= 12'h555;
      20'h075f5: out <= 12'h555;
      20'h075f6: out <= 12'h555;
      20'h075f7: out <= 12'h555;
      20'h075f8: out <= 12'h555;
      20'h075f9: out <= 12'h555;
      20'h075fa: out <= 12'h555;
      20'h075fb: out <= 12'h555;
      20'h075fc: out <= 12'h555;
      20'h075fd: out <= 12'h555;
      20'h075fe: out <= 12'h555;
      20'h075ff: out <= 12'h777;
      20'h07600: out <= 12'h000;
      20'h07601: out <= 12'h000;
      20'h07602: out <= 12'h000;
      20'h07603: out <= 12'h000;
      20'h07604: out <= 12'hf87;
      20'h07605: out <= 12'h000;
      20'h07606: out <= 12'h000;
      20'h07607: out <= 12'h000;
      20'h07608: out <= 12'hfa9;
      20'h07609: out <= 12'hfa9;
      20'h0760a: out <= 12'hfa9;
      20'h0760b: out <= 12'hfa9;
      20'h0760c: out <= 12'hfa9;
      20'h0760d: out <= 12'hfa9;
      20'h0760e: out <= 12'hfa9;
      20'h0760f: out <= 12'hfa9;
      20'h07610: out <= 12'hf76;
      20'h07611: out <= 12'hf76;
      20'h07612: out <= 12'hf76;
      20'h07613: out <= 12'hf76;
      20'h07614: out <= 12'hf76;
      20'h07615: out <= 12'hf76;
      20'h07616: out <= 12'hf76;
      20'h07617: out <= 12'hf76;
      20'h07618: out <= 12'h000;
      20'h07619: out <= 12'h000;
      20'h0761a: out <= 12'h000;
      20'h0761b: out <= 12'h000;
      20'h0761c: out <= 12'h000;
      20'h0761d: out <= 12'h000;
      20'h0761e: out <= 12'h000;
      20'h0761f: out <= 12'h000;
      20'h07620: out <= 12'h222;
      20'h07621: out <= 12'h222;
      20'h07622: out <= 12'hbbb;
      20'h07623: out <= 12'h666;
      20'h07624: out <= 12'hbbb;
      20'h07625: out <= 12'h666;
      20'h07626: out <= 12'hbbb;
      20'h07627: out <= 12'h666;
      20'h07628: out <= 12'hbbb;
      20'h07629: out <= 12'h666;
      20'h0762a: out <= 12'hbbb;
      20'h0762b: out <= 12'h666;
      20'h0762c: out <= 12'hbbb;
      20'h0762d: out <= 12'h222;
      20'h0762e: out <= 12'h222;
      20'h0762f: out <= 12'h222;
      20'h07630: out <= 12'h000;
      20'h07631: out <= 12'h000;
      20'h07632: out <= 12'h666;
      20'h07633: out <= 12'hbbb;
      20'h07634: out <= 12'h666;
      20'h07635: out <= 12'hbbb;
      20'h07636: out <= 12'h666;
      20'h07637: out <= 12'hbbb;
      20'h07638: out <= 12'h666;
      20'h07639: out <= 12'hbbb;
      20'h0763a: out <= 12'h666;
      20'h0763b: out <= 12'hbbb;
      20'h0763c: out <= 12'h666;
      20'h0763d: out <= 12'h000;
      20'h0763e: out <= 12'h000;
      20'h0763f: out <= 12'h000;
      20'h07640: out <= 12'h222;
      20'h07641: out <= 12'h222;
      20'h07642: out <= 12'h666;
      20'h07643: out <= 12'h666;
      20'h07644: out <= 12'h666;
      20'h07645: out <= 12'hfff;
      20'h07646: out <= 12'hfff;
      20'h07647: out <= 12'hbbb;
      20'h07648: out <= 12'hbbb;
      20'h07649: out <= 12'hbbb;
      20'h0764a: out <= 12'h666;
      20'h0764b: out <= 12'h666;
      20'h0764c: out <= 12'h666;
      20'h0764d: out <= 12'h666;
      20'h0764e: out <= 12'h666;
      20'h0764f: out <= 12'h222;
      20'h07650: out <= 12'h000;
      20'h07651: out <= 12'h000;
      20'h07652: out <= 12'h666;
      20'h07653: out <= 12'hbbb;
      20'h07654: out <= 12'h666;
      20'h07655: out <= 12'hfff;
      20'h07656: out <= 12'hfff;
      20'h07657: out <= 12'hbbb;
      20'h07658: out <= 12'hbbb;
      20'h07659: out <= 12'hbbb;
      20'h0765a: out <= 12'h666;
      20'h0765b: out <= 12'h666;
      20'h0765c: out <= 12'h666;
      20'h0765d: out <= 12'hbbb;
      20'h0765e: out <= 12'h666;
      20'h0765f: out <= 12'h000;
      20'h07660: out <= 12'h222;
      20'h07661: out <= 12'h222;
      20'h07662: out <= 12'h222;
      20'h07663: out <= 12'hbbb;
      20'h07664: out <= 12'h666;
      20'h07665: out <= 12'hbbb;
      20'h07666: out <= 12'h666;
      20'h07667: out <= 12'hbbb;
      20'h07668: out <= 12'h666;
      20'h07669: out <= 12'hbbb;
      20'h0766a: out <= 12'h666;
      20'h0766b: out <= 12'hbbb;
      20'h0766c: out <= 12'h666;
      20'h0766d: out <= 12'hbbb;
      20'h0766e: out <= 12'h222;
      20'h0766f: out <= 12'h222;
      20'h07670: out <= 12'h000;
      20'h07671: out <= 12'h000;
      20'h07672: out <= 12'h000;
      20'h07673: out <= 12'h666;
      20'h07674: out <= 12'hbbb;
      20'h07675: out <= 12'h666;
      20'h07676: out <= 12'hbbb;
      20'h07677: out <= 12'h666;
      20'h07678: out <= 12'hbbb;
      20'h07679: out <= 12'h666;
      20'h0767a: out <= 12'hbbb;
      20'h0767b: out <= 12'h666;
      20'h0767c: out <= 12'hbbb;
      20'h0767d: out <= 12'h666;
      20'h0767e: out <= 12'h000;
      20'h0767f: out <= 12'h000;
      20'h07680: out <= 12'h222;
      20'h07681: out <= 12'h222;
      20'h07682: out <= 12'h222;
      20'h07683: out <= 12'hbbb;
      20'h07684: out <= 12'h222;
      20'h07685: out <= 12'h666;
      20'h07686: out <= 12'h666;
      20'h07687: out <= 12'hbbb;
      20'h07688: out <= 12'hfff;
      20'h07689: out <= 12'hbbb;
      20'h0768a: out <= 12'h666;
      20'h0768b: out <= 12'h666;
      20'h0768c: out <= 12'h222;
      20'h0768d: out <= 12'hbbb;
      20'h0768e: out <= 12'h222;
      20'h0768f: out <= 12'h222;
      20'h07690: out <= 12'h000;
      20'h07691: out <= 12'h000;
      20'h07692: out <= 12'h000;
      20'h07693: out <= 12'h666;
      20'h07694: out <= 12'h000;
      20'h07695: out <= 12'h666;
      20'h07696: out <= 12'h666;
      20'h07697: out <= 12'hbbb;
      20'h07698: out <= 12'hfff;
      20'h07699: out <= 12'hbbb;
      20'h0769a: out <= 12'h666;
      20'h0769b: out <= 12'h666;
      20'h0769c: out <= 12'h000;
      20'h0769d: out <= 12'h666;
      20'h0769e: out <= 12'h000;
      20'h0769f: out <= 12'h000;
      20'h076a0: out <= 12'h603;
      20'h076a1: out <= 12'h603;
      20'h076a2: out <= 12'h603;
      20'h076a3: out <= 12'h603;
      20'h076a4: out <= 12'h603;
      20'h076a5: out <= 12'h603;
      20'h076a6: out <= 12'h603;
      20'h076a7: out <= 12'h603;
      20'h076a8: out <= 12'h603;
      20'h076a9: out <= 12'h603;
      20'h076aa: out <= 12'h603;
      20'h076ab: out <= 12'h603;
      20'h076ac: out <= 12'hee9;
      20'h076ad: out <= 12'hf87;
      20'h076ae: out <= 12'hee9;
      20'h076af: out <= 12'hf87;
      20'h076b0: out <= 12'hf87;
      20'h076b1: out <= 12'hb27;
      20'h076b2: out <= 12'hf87;
      20'h076b3: out <= 12'hb27;
      20'h076b4: out <= 12'h603;
      20'h076b5: out <= 12'h603;
      20'h076b6: out <= 12'h603;
      20'h076b7: out <= 12'h603;
      20'h076b8: out <= 12'h603;
      20'h076b9: out <= 12'h603;
      20'h076ba: out <= 12'h603;
      20'h076bb: out <= 12'h603;
      20'h076bc: out <= 12'h603;
      20'h076bd: out <= 12'h603;
      20'h076be: out <= 12'h603;
      20'h076bf: out <= 12'h603;
      20'h076c0: out <= 12'h603;
      20'h076c1: out <= 12'h603;
      20'h076c2: out <= 12'h603;
      20'h076c3: out <= 12'h603;
      20'h076c4: out <= 12'hee9;
      20'h076c5: out <= 12'hf87;
      20'h076c6: out <= 12'hee9;
      20'h076c7: out <= 12'hf87;
      20'h076c8: out <= 12'hf87;
      20'h076c9: out <= 12'hb27;
      20'h076ca: out <= 12'hf87;
      20'h076cb: out <= 12'hb27;
      20'h076cc: out <= 12'h603;
      20'h076cd: out <= 12'h603;
      20'h076ce: out <= 12'h603;
      20'h076cf: out <= 12'h603;
      20'h076d0: out <= 12'h603;
      20'h076d1: out <= 12'h603;
      20'h076d2: out <= 12'h603;
      20'h076d3: out <= 12'h603;
      20'h076d4: out <= 12'h603;
      20'h076d5: out <= 12'h603;
      20'h076d6: out <= 12'h603;
      20'h076d7: out <= 12'h603;
      20'h076d8: out <= 12'h603;
      20'h076d9: out <= 12'h603;
      20'h076da: out <= 12'h603;
      20'h076db: out <= 12'h603;
      20'h076dc: out <= 12'h603;
      20'h076dd: out <= 12'h603;
      20'h076de: out <= 12'h603;
      20'h076df: out <= 12'h603;
      20'h076e0: out <= 12'h603;
      20'h076e1: out <= 12'h603;
      20'h076e2: out <= 12'h603;
      20'h076e3: out <= 12'h603;
      20'h076e4: out <= 12'h603;
      20'h076e5: out <= 12'h603;
      20'h076e6: out <= 12'h603;
      20'h076e7: out <= 12'h603;
      20'h076e8: out <= 12'h603;
      20'h076e9: out <= 12'h603;
      20'h076ea: out <= 12'h603;
      20'h076eb: out <= 12'h603;
      20'h076ec: out <= 12'h603;
      20'h076ed: out <= 12'h603;
      20'h076ee: out <= 12'h603;
      20'h076ef: out <= 12'h603;
      20'h076f0: out <= 12'h603;
      20'h076f1: out <= 12'h603;
      20'h076f2: out <= 12'h603;
      20'h076f3: out <= 12'h603;
      20'h076f4: out <= 12'h603;
      20'h076f5: out <= 12'h603;
      20'h076f6: out <= 12'h603;
      20'h076f7: out <= 12'h603;
      20'h076f8: out <= 12'hee9;
      20'h076f9: out <= 12'hf87;
      20'h076fa: out <= 12'hee9;
      20'h076fb: out <= 12'hf87;
      20'h076fc: out <= 12'hf87;
      20'h076fd: out <= 12'hb27;
      20'h076fe: out <= 12'hf87;
      20'h076ff: out <= 12'hb27;
      20'h07700: out <= 12'h000;
      20'h07701: out <= 12'h000;
      20'h07702: out <= 12'h000;
      20'h07703: out <= 12'h000;
      20'h07704: out <= 12'h000;
      20'h07705: out <= 12'h000;
      20'h07706: out <= 12'h000;
      20'h07707: out <= 12'h000;
      20'h07708: out <= 12'h777;
      20'h07709: out <= 12'h555;
      20'h0770a: out <= 12'h555;
      20'h0770b: out <= 12'h555;
      20'h0770c: out <= 12'h555;
      20'h0770d: out <= 12'h555;
      20'h0770e: out <= 12'h555;
      20'h0770f: out <= 12'h555;
      20'h07710: out <= 12'h555;
      20'h07711: out <= 12'h555;
      20'h07712: out <= 12'h555;
      20'h07713: out <= 12'h555;
      20'h07714: out <= 12'h555;
      20'h07715: out <= 12'h555;
      20'h07716: out <= 12'h555;
      20'h07717: out <= 12'h777;
      20'h07718: out <= 12'h000;
      20'h07719: out <= 12'h000;
      20'h0771a: out <= 12'h000;
      20'h0771b: out <= 12'hf87;
      20'h0771c: out <= 12'h000;
      20'h0771d: out <= 12'hf87;
      20'h0771e: out <= 12'h000;
      20'h0771f: out <= 12'h000;
      20'h07720: out <= 12'hfa9;
      20'h07721: out <= 12'hfa9;
      20'h07722: out <= 12'hfa9;
      20'h07723: out <= 12'hfa9;
      20'h07724: out <= 12'hfa9;
      20'h07725: out <= 12'hfa9;
      20'h07726: out <= 12'hfa9;
      20'h07727: out <= 12'hfa9;
      20'h07728: out <= 12'hf76;
      20'h07729: out <= 12'hf76;
      20'h0772a: out <= 12'hf76;
      20'h0772b: out <= 12'hf76;
      20'h0772c: out <= 12'hf76;
      20'h0772d: out <= 12'hf76;
      20'h0772e: out <= 12'hf76;
      20'h0772f: out <= 12'hf76;
      20'h07730: out <= 12'h000;
      20'h07731: out <= 12'h000;
      20'h07732: out <= 12'h000;
      20'h07733: out <= 12'h000;
      20'h07734: out <= 12'h000;
      20'h07735: out <= 12'h000;
      20'h07736: out <= 12'h000;
      20'h07737: out <= 12'h000;
      20'h07738: out <= 12'h222;
      20'h07739: out <= 12'h222;
      20'h0773a: out <= 12'h222;
      20'h0773b: out <= 12'h666;
      20'h0773c: out <= 12'h222;
      20'h0773d: out <= 12'h666;
      20'h0773e: out <= 12'h222;
      20'h0773f: out <= 12'h666;
      20'h07740: out <= 12'h222;
      20'h07741: out <= 12'h666;
      20'h07742: out <= 12'h222;
      20'h07743: out <= 12'h666;
      20'h07744: out <= 12'h222;
      20'h07745: out <= 12'h222;
      20'h07746: out <= 12'h222;
      20'h07747: out <= 12'h222;
      20'h07748: out <= 12'h000;
      20'h07749: out <= 12'h000;
      20'h0774a: out <= 12'h000;
      20'h0774b: out <= 12'h666;
      20'h0774c: out <= 12'h000;
      20'h0774d: out <= 12'h666;
      20'h0774e: out <= 12'h000;
      20'h0774f: out <= 12'h666;
      20'h07750: out <= 12'h000;
      20'h07751: out <= 12'h666;
      20'h07752: out <= 12'h000;
      20'h07753: out <= 12'h666;
      20'h07754: out <= 12'h000;
      20'h07755: out <= 12'h000;
      20'h07756: out <= 12'h000;
      20'h07757: out <= 12'h000;
      20'h07758: out <= 12'h222;
      20'h07759: out <= 12'h222;
      20'h0775a: out <= 12'h222;
      20'h0775b: out <= 12'hbbb;
      20'h0775c: out <= 12'h222;
      20'h0775d: out <= 12'h666;
      20'h0775e: out <= 12'hfff;
      20'h0775f: out <= 12'hbbb;
      20'h07760: out <= 12'hbbb;
      20'h07761: out <= 12'hbbb;
      20'h07762: out <= 12'h666;
      20'h07763: out <= 12'h666;
      20'h07764: out <= 12'h222;
      20'h07765: out <= 12'hbbb;
      20'h07766: out <= 12'h222;
      20'h07767: out <= 12'h222;
      20'h07768: out <= 12'h000;
      20'h07769: out <= 12'h000;
      20'h0776a: out <= 12'h000;
      20'h0776b: out <= 12'h666;
      20'h0776c: out <= 12'h000;
      20'h0776d: out <= 12'h666;
      20'h0776e: out <= 12'hfff;
      20'h0776f: out <= 12'hbbb;
      20'h07770: out <= 12'hbbb;
      20'h07771: out <= 12'hbbb;
      20'h07772: out <= 12'h666;
      20'h07773: out <= 12'h666;
      20'h07774: out <= 12'h000;
      20'h07775: out <= 12'h666;
      20'h07776: out <= 12'h000;
      20'h07777: out <= 12'h000;
      20'h07778: out <= 12'h222;
      20'h07779: out <= 12'h222;
      20'h0777a: out <= 12'h222;
      20'h0777b: out <= 12'h222;
      20'h0777c: out <= 12'h666;
      20'h0777d: out <= 12'h222;
      20'h0777e: out <= 12'h666;
      20'h0777f: out <= 12'h222;
      20'h07780: out <= 12'h666;
      20'h07781: out <= 12'h222;
      20'h07782: out <= 12'h666;
      20'h07783: out <= 12'h222;
      20'h07784: out <= 12'h666;
      20'h07785: out <= 12'h222;
      20'h07786: out <= 12'h222;
      20'h07787: out <= 12'h222;
      20'h07788: out <= 12'h000;
      20'h07789: out <= 12'h000;
      20'h0778a: out <= 12'h000;
      20'h0778b: out <= 12'h000;
      20'h0778c: out <= 12'h666;
      20'h0778d: out <= 12'h000;
      20'h0778e: out <= 12'h666;
      20'h0778f: out <= 12'h000;
      20'h07790: out <= 12'h666;
      20'h07791: out <= 12'h000;
      20'h07792: out <= 12'h666;
      20'h07793: out <= 12'h000;
      20'h07794: out <= 12'h666;
      20'h07795: out <= 12'h000;
      20'h07796: out <= 12'h000;
      20'h07797: out <= 12'h000;
      20'h07798: out <= 12'h222;
      20'h07799: out <= 12'h222;
      20'h0779a: out <= 12'h222;
      20'h0779b: out <= 12'h222;
      20'h0779c: out <= 12'h222;
      20'h0779d: out <= 12'h222;
      20'h0779e: out <= 12'h666;
      20'h0779f: out <= 12'hbbb;
      20'h077a0: out <= 12'hfff;
      20'h077a1: out <= 12'hbbb;
      20'h077a2: out <= 12'h666;
      20'h077a3: out <= 12'h222;
      20'h077a4: out <= 12'h222;
      20'h077a5: out <= 12'h222;
      20'h077a6: out <= 12'h222;
      20'h077a7: out <= 12'h222;
      20'h077a8: out <= 12'h000;
      20'h077a9: out <= 12'h000;
      20'h077aa: out <= 12'h000;
      20'h077ab: out <= 12'h000;
      20'h077ac: out <= 12'h000;
      20'h077ad: out <= 12'h000;
      20'h077ae: out <= 12'h666;
      20'h077af: out <= 12'hbbb;
      20'h077b0: out <= 12'hfff;
      20'h077b1: out <= 12'hbbb;
      20'h077b2: out <= 12'h666;
      20'h077b3: out <= 12'h000;
      20'h077b4: out <= 12'h000;
      20'h077b5: out <= 12'h000;
      20'h077b6: out <= 12'h000;
      20'h077b7: out <= 12'h000;
      20'h077b8: out <= 12'h603;
      20'h077b9: out <= 12'h603;
      20'h077ba: out <= 12'h603;
      20'h077bb: out <= 12'h603;
      20'h077bc: out <= 12'h603;
      20'h077bd: out <= 12'h603;
      20'h077be: out <= 12'h603;
      20'h077bf: out <= 12'h603;
      20'h077c0: out <= 12'h603;
      20'h077c1: out <= 12'h603;
      20'h077c2: out <= 12'h603;
      20'h077c3: out <= 12'h603;
      20'h077c4: out <= 12'hee9;
      20'h077c5: out <= 12'hf87;
      20'h077c6: out <= 12'hee9;
      20'h077c7: out <= 12'hb27;
      20'h077c8: out <= 12'hb27;
      20'h077c9: out <= 12'hb27;
      20'h077ca: out <= 12'hf87;
      20'h077cb: out <= 12'hb27;
      20'h077cc: out <= 12'h603;
      20'h077cd: out <= 12'h603;
      20'h077ce: out <= 12'h603;
      20'h077cf: out <= 12'h603;
      20'h077d0: out <= 12'h603;
      20'h077d1: out <= 12'h603;
      20'h077d2: out <= 12'h603;
      20'h077d3: out <= 12'h603;
      20'h077d4: out <= 12'h603;
      20'h077d5: out <= 12'h603;
      20'h077d6: out <= 12'h603;
      20'h077d7: out <= 12'h603;
      20'h077d8: out <= 12'h603;
      20'h077d9: out <= 12'h603;
      20'h077da: out <= 12'h603;
      20'h077db: out <= 12'h603;
      20'h077dc: out <= 12'hee9;
      20'h077dd: out <= 12'hf87;
      20'h077de: out <= 12'hee9;
      20'h077df: out <= 12'hb27;
      20'h077e0: out <= 12'hb27;
      20'h077e1: out <= 12'hb27;
      20'h077e2: out <= 12'hf87;
      20'h077e3: out <= 12'hb27;
      20'h077e4: out <= 12'h603;
      20'h077e5: out <= 12'h603;
      20'h077e6: out <= 12'h603;
      20'h077e7: out <= 12'h603;
      20'h077e8: out <= 12'h603;
      20'h077e9: out <= 12'h603;
      20'h077ea: out <= 12'h603;
      20'h077eb: out <= 12'h603;
      20'h077ec: out <= 12'h603;
      20'h077ed: out <= 12'h603;
      20'h077ee: out <= 12'h603;
      20'h077ef: out <= 12'h603;
      20'h077f0: out <= 12'h603;
      20'h077f1: out <= 12'h603;
      20'h077f2: out <= 12'h603;
      20'h077f3: out <= 12'h603;
      20'h077f4: out <= 12'h603;
      20'h077f5: out <= 12'h603;
      20'h077f6: out <= 12'h603;
      20'h077f7: out <= 12'h603;
      20'h077f8: out <= 12'h603;
      20'h077f9: out <= 12'h603;
      20'h077fa: out <= 12'h603;
      20'h077fb: out <= 12'h603;
      20'h077fc: out <= 12'h603;
      20'h077fd: out <= 12'h603;
      20'h077fe: out <= 12'h603;
      20'h077ff: out <= 12'h603;
      20'h07800: out <= 12'h603;
      20'h07801: out <= 12'h603;
      20'h07802: out <= 12'h603;
      20'h07803: out <= 12'h603;
      20'h07804: out <= 12'h603;
      20'h07805: out <= 12'h603;
      20'h07806: out <= 12'h603;
      20'h07807: out <= 12'h603;
      20'h07808: out <= 12'h603;
      20'h07809: out <= 12'h603;
      20'h0780a: out <= 12'h603;
      20'h0780b: out <= 12'h603;
      20'h0780c: out <= 12'h603;
      20'h0780d: out <= 12'h603;
      20'h0780e: out <= 12'h603;
      20'h0780f: out <= 12'h603;
      20'h07810: out <= 12'hee9;
      20'h07811: out <= 12'hf87;
      20'h07812: out <= 12'hee9;
      20'h07813: out <= 12'hb27;
      20'h07814: out <= 12'hb27;
      20'h07815: out <= 12'hb27;
      20'h07816: out <= 12'hf87;
      20'h07817: out <= 12'hb27;
      20'h07818: out <= 12'h000;
      20'h07819: out <= 12'h000;
      20'h0781a: out <= 12'h000;
      20'h0781b: out <= 12'h000;
      20'h0781c: out <= 12'h000;
      20'h0781d: out <= 12'h000;
      20'h0781e: out <= 12'h000;
      20'h0781f: out <= 12'h000;
      20'h07820: out <= 12'h777;
      20'h07821: out <= 12'h555;
      20'h07822: out <= 12'h555;
      20'h07823: out <= 12'h555;
      20'h07824: out <= 12'h555;
      20'h07825: out <= 12'h555;
      20'h07826: out <= 12'h555;
      20'h07827: out <= 12'h555;
      20'h07828: out <= 12'h555;
      20'h07829: out <= 12'h555;
      20'h0782a: out <= 12'h555;
      20'h0782b: out <= 12'h555;
      20'h0782c: out <= 12'h555;
      20'h0782d: out <= 12'h555;
      20'h0782e: out <= 12'h555;
      20'h0782f: out <= 12'h777;
      20'h07830: out <= 12'h000;
      20'h07831: out <= 12'h000;
      20'h07832: out <= 12'hf87;
      20'h07833: out <= 12'h000;
      20'h07834: out <= 12'h000;
      20'h07835: out <= 12'h000;
      20'h07836: out <= 12'hf87;
      20'h07837: out <= 12'h000;
      20'h07838: out <= 12'hfa9;
      20'h07839: out <= 12'hfa9;
      20'h0783a: out <= 12'hfa9;
      20'h0783b: out <= 12'hfa9;
      20'h0783c: out <= 12'hfa9;
      20'h0783d: out <= 12'hfa9;
      20'h0783e: out <= 12'hfa9;
      20'h0783f: out <= 12'hfa9;
      20'h07840: out <= 12'hf76;
      20'h07841: out <= 12'hf76;
      20'h07842: out <= 12'hf76;
      20'h07843: out <= 12'hf76;
      20'h07844: out <= 12'hf76;
      20'h07845: out <= 12'hf76;
      20'h07846: out <= 12'hf76;
      20'h07847: out <= 12'hf76;
      20'h07848: out <= 12'h000;
      20'h07849: out <= 12'h000;
      20'h0784a: out <= 12'h000;
      20'h0784b: out <= 12'h000;
      20'h0784c: out <= 12'h000;
      20'h0784d: out <= 12'h000;
      20'h0784e: out <= 12'h000;
      20'h0784f: out <= 12'h000;
      20'h07850: out <= 12'h222;
      20'h07851: out <= 12'h222;
      20'h07852: out <= 12'h222;
      20'h07853: out <= 12'h222;
      20'h07854: out <= 12'h222;
      20'h07855: out <= 12'h222;
      20'h07856: out <= 12'h222;
      20'h07857: out <= 12'h222;
      20'h07858: out <= 12'h222;
      20'h07859: out <= 12'h222;
      20'h0785a: out <= 12'h222;
      20'h0785b: out <= 12'h222;
      20'h0785c: out <= 12'h222;
      20'h0785d: out <= 12'h222;
      20'h0785e: out <= 12'h222;
      20'h0785f: out <= 12'h222;
      20'h07860: out <= 12'h000;
      20'h07861: out <= 12'h000;
      20'h07862: out <= 12'h000;
      20'h07863: out <= 12'h000;
      20'h07864: out <= 12'h000;
      20'h07865: out <= 12'h000;
      20'h07866: out <= 12'h000;
      20'h07867: out <= 12'h000;
      20'h07868: out <= 12'h000;
      20'h07869: out <= 12'h000;
      20'h0786a: out <= 12'h000;
      20'h0786b: out <= 12'h000;
      20'h0786c: out <= 12'h000;
      20'h0786d: out <= 12'h000;
      20'h0786e: out <= 12'h000;
      20'h0786f: out <= 12'h000;
      20'h07870: out <= 12'h222;
      20'h07871: out <= 12'h222;
      20'h07872: out <= 12'h222;
      20'h07873: out <= 12'h222;
      20'h07874: out <= 12'h222;
      20'h07875: out <= 12'h222;
      20'h07876: out <= 12'h666;
      20'h07877: out <= 12'h666;
      20'h07878: out <= 12'h666;
      20'h07879: out <= 12'h666;
      20'h0787a: out <= 12'h666;
      20'h0787b: out <= 12'h222;
      20'h0787c: out <= 12'h222;
      20'h0787d: out <= 12'h222;
      20'h0787e: out <= 12'h222;
      20'h0787f: out <= 12'h222;
      20'h07880: out <= 12'h000;
      20'h07881: out <= 12'h000;
      20'h07882: out <= 12'h000;
      20'h07883: out <= 12'h000;
      20'h07884: out <= 12'h000;
      20'h07885: out <= 12'h000;
      20'h07886: out <= 12'h666;
      20'h07887: out <= 12'h666;
      20'h07888: out <= 12'h666;
      20'h07889: out <= 12'h666;
      20'h0788a: out <= 12'h666;
      20'h0788b: out <= 12'h000;
      20'h0788c: out <= 12'h000;
      20'h0788d: out <= 12'h000;
      20'h0788e: out <= 12'h000;
      20'h0788f: out <= 12'h000;
      20'h07890: out <= 12'h222;
      20'h07891: out <= 12'h222;
      20'h07892: out <= 12'h222;
      20'h07893: out <= 12'h222;
      20'h07894: out <= 12'h222;
      20'h07895: out <= 12'h222;
      20'h07896: out <= 12'h222;
      20'h07897: out <= 12'h222;
      20'h07898: out <= 12'h222;
      20'h07899: out <= 12'h222;
      20'h0789a: out <= 12'h222;
      20'h0789b: out <= 12'h222;
      20'h0789c: out <= 12'h222;
      20'h0789d: out <= 12'h222;
      20'h0789e: out <= 12'h222;
      20'h0789f: out <= 12'h222;
      20'h078a0: out <= 12'h000;
      20'h078a1: out <= 12'h000;
      20'h078a2: out <= 12'h000;
      20'h078a3: out <= 12'h000;
      20'h078a4: out <= 12'h000;
      20'h078a5: out <= 12'h000;
      20'h078a6: out <= 12'h000;
      20'h078a7: out <= 12'h000;
      20'h078a8: out <= 12'h000;
      20'h078a9: out <= 12'h000;
      20'h078aa: out <= 12'h000;
      20'h078ab: out <= 12'h000;
      20'h078ac: out <= 12'h000;
      20'h078ad: out <= 12'h000;
      20'h078ae: out <= 12'h000;
      20'h078af: out <= 12'h000;
      20'h078b0: out <= 12'h222;
      20'h078b1: out <= 12'h222;
      20'h078b2: out <= 12'h222;
      20'h078b3: out <= 12'h222;
      20'h078b4: out <= 12'h222;
      20'h078b5: out <= 12'h222;
      20'h078b6: out <= 12'h666;
      20'h078b7: out <= 12'hbbb;
      20'h078b8: out <= 12'hfff;
      20'h078b9: out <= 12'hbbb;
      20'h078ba: out <= 12'h666;
      20'h078bb: out <= 12'h222;
      20'h078bc: out <= 12'h222;
      20'h078bd: out <= 12'h222;
      20'h078be: out <= 12'h222;
      20'h078bf: out <= 12'h222;
      20'h078c0: out <= 12'h000;
      20'h078c1: out <= 12'h000;
      20'h078c2: out <= 12'h000;
      20'h078c3: out <= 12'h000;
      20'h078c4: out <= 12'h000;
      20'h078c5: out <= 12'h000;
      20'h078c6: out <= 12'h666;
      20'h078c7: out <= 12'hbbb;
      20'h078c8: out <= 12'hfff;
      20'h078c9: out <= 12'hbbb;
      20'h078ca: out <= 12'h666;
      20'h078cb: out <= 12'h000;
      20'h078cc: out <= 12'h000;
      20'h078cd: out <= 12'h000;
      20'h078ce: out <= 12'h000;
      20'h078cf: out <= 12'h000;
      20'h078d0: out <= 12'h603;
      20'h078d1: out <= 12'h603;
      20'h078d2: out <= 12'h603;
      20'h078d3: out <= 12'h603;
      20'h078d4: out <= 12'h603;
      20'h078d5: out <= 12'h603;
      20'h078d6: out <= 12'h603;
      20'h078d7: out <= 12'h603;
      20'h078d8: out <= 12'h603;
      20'h078d9: out <= 12'h603;
      20'h078da: out <= 12'h603;
      20'h078db: out <= 12'h603;
      20'h078dc: out <= 12'hee9;
      20'h078dd: out <= 12'hf87;
      20'h078de: out <= 12'hf87;
      20'h078df: out <= 12'hf87;
      20'h078e0: out <= 12'hf87;
      20'h078e1: out <= 12'hf87;
      20'h078e2: out <= 12'hf87;
      20'h078e3: out <= 12'hb27;
      20'h078e4: out <= 12'h603;
      20'h078e5: out <= 12'h603;
      20'h078e6: out <= 12'h603;
      20'h078e7: out <= 12'h603;
      20'h078e8: out <= 12'h603;
      20'h078e9: out <= 12'h603;
      20'h078ea: out <= 12'h603;
      20'h078eb: out <= 12'h603;
      20'h078ec: out <= 12'h603;
      20'h078ed: out <= 12'h603;
      20'h078ee: out <= 12'h603;
      20'h078ef: out <= 12'h603;
      20'h078f0: out <= 12'h603;
      20'h078f1: out <= 12'h603;
      20'h078f2: out <= 12'h603;
      20'h078f3: out <= 12'h603;
      20'h078f4: out <= 12'hee9;
      20'h078f5: out <= 12'hf87;
      20'h078f6: out <= 12'hf87;
      20'h078f7: out <= 12'hf87;
      20'h078f8: out <= 12'hf87;
      20'h078f9: out <= 12'hf87;
      20'h078fa: out <= 12'hf87;
      20'h078fb: out <= 12'hb27;
      20'h078fc: out <= 12'h603;
      20'h078fd: out <= 12'h603;
      20'h078fe: out <= 12'h603;
      20'h078ff: out <= 12'h603;
      20'h07900: out <= 12'h603;
      20'h07901: out <= 12'h603;
      20'h07902: out <= 12'h603;
      20'h07903: out <= 12'h603;
      20'h07904: out <= 12'h603;
      20'h07905: out <= 12'h603;
      20'h07906: out <= 12'h603;
      20'h07907: out <= 12'h603;
      20'h07908: out <= 12'h603;
      20'h07909: out <= 12'h603;
      20'h0790a: out <= 12'h603;
      20'h0790b: out <= 12'h603;
      20'h0790c: out <= 12'h603;
      20'h0790d: out <= 12'h603;
      20'h0790e: out <= 12'h603;
      20'h0790f: out <= 12'h603;
      20'h07910: out <= 12'h603;
      20'h07911: out <= 12'h603;
      20'h07912: out <= 12'h603;
      20'h07913: out <= 12'h603;
      20'h07914: out <= 12'h603;
      20'h07915: out <= 12'h603;
      20'h07916: out <= 12'h603;
      20'h07917: out <= 12'h603;
      20'h07918: out <= 12'h603;
      20'h07919: out <= 12'h603;
      20'h0791a: out <= 12'h603;
      20'h0791b: out <= 12'h603;
      20'h0791c: out <= 12'h603;
      20'h0791d: out <= 12'h603;
      20'h0791e: out <= 12'h603;
      20'h0791f: out <= 12'h603;
      20'h07920: out <= 12'h603;
      20'h07921: out <= 12'h603;
      20'h07922: out <= 12'h603;
      20'h07923: out <= 12'h603;
      20'h07924: out <= 12'h603;
      20'h07925: out <= 12'h603;
      20'h07926: out <= 12'h603;
      20'h07927: out <= 12'h603;
      20'h07928: out <= 12'hee9;
      20'h07929: out <= 12'hf87;
      20'h0792a: out <= 12'hf87;
      20'h0792b: out <= 12'hf87;
      20'h0792c: out <= 12'hf87;
      20'h0792d: out <= 12'hf87;
      20'h0792e: out <= 12'hf87;
      20'h0792f: out <= 12'hb27;
      20'h07930: out <= 12'h000;
      20'h07931: out <= 12'h000;
      20'h07932: out <= 12'h000;
      20'h07933: out <= 12'h000;
      20'h07934: out <= 12'h000;
      20'h07935: out <= 12'h000;
      20'h07936: out <= 12'h000;
      20'h07937: out <= 12'h000;
      20'h07938: out <= 12'h777;
      20'h07939: out <= 12'h777;
      20'h0793a: out <= 12'h555;
      20'h0793b: out <= 12'h555;
      20'h0793c: out <= 12'h555;
      20'h0793d: out <= 12'h555;
      20'h0793e: out <= 12'h555;
      20'h0793f: out <= 12'h555;
      20'h07940: out <= 12'h555;
      20'h07941: out <= 12'h555;
      20'h07942: out <= 12'h555;
      20'h07943: out <= 12'h555;
      20'h07944: out <= 12'h555;
      20'h07945: out <= 12'h555;
      20'h07946: out <= 12'h777;
      20'h07947: out <= 12'h777;
      20'h07948: out <= 12'h000;
      20'h07949: out <= 12'h000;
      20'h0794a: out <= 12'h000;
      20'h0794b: out <= 12'h000;
      20'h0794c: out <= 12'h000;
      20'h0794d: out <= 12'h000;
      20'h0794e: out <= 12'h000;
      20'h0794f: out <= 12'h000;
      20'h07950: out <= 12'hfa9;
      20'h07951: out <= 12'hfa9;
      20'h07952: out <= 12'hfa9;
      20'h07953: out <= 12'hfa9;
      20'h07954: out <= 12'hfa9;
      20'h07955: out <= 12'hfa9;
      20'h07956: out <= 12'hfa9;
      20'h07957: out <= 12'hfa9;
      20'h07958: out <= 12'hf76;
      20'h07959: out <= 12'hf76;
      20'h0795a: out <= 12'hf76;
      20'h0795b: out <= 12'hf76;
      20'h0795c: out <= 12'hf76;
      20'h0795d: out <= 12'hf76;
      20'h0795e: out <= 12'hf76;
      20'h0795f: out <= 12'hf76;
      20'h07960: out <= 12'h000;
      20'h07961: out <= 12'h000;
      20'h07962: out <= 12'h000;
      20'h07963: out <= 12'h000;
      20'h07964: out <= 12'h000;
      20'h07965: out <= 12'h000;
      20'h07966: out <= 12'h000;
      20'h07967: out <= 12'h000;
      20'h07968: out <= 12'h222;
      20'h07969: out <= 12'h222;
      20'h0796a: out <= 12'h222;
      20'h0796b: out <= 12'h222;
      20'h0796c: out <= 12'h222;
      20'h0796d: out <= 12'h222;
      20'h0796e: out <= 12'h222;
      20'h0796f: out <= 12'h222;
      20'h07970: out <= 12'h222;
      20'h07971: out <= 12'h222;
      20'h07972: out <= 12'h222;
      20'h07973: out <= 12'h222;
      20'h07974: out <= 12'h222;
      20'h07975: out <= 12'h222;
      20'h07976: out <= 12'h222;
      20'h07977: out <= 12'h222;
      20'h07978: out <= 12'h000;
      20'h07979: out <= 12'h000;
      20'h0797a: out <= 12'h000;
      20'h0797b: out <= 12'h000;
      20'h0797c: out <= 12'h000;
      20'h0797d: out <= 12'h000;
      20'h0797e: out <= 12'h000;
      20'h0797f: out <= 12'h000;
      20'h07980: out <= 12'h000;
      20'h07981: out <= 12'h000;
      20'h07982: out <= 12'h000;
      20'h07983: out <= 12'h000;
      20'h07984: out <= 12'h000;
      20'h07985: out <= 12'h000;
      20'h07986: out <= 12'h000;
      20'h07987: out <= 12'h000;
      20'h07988: out <= 12'h222;
      20'h07989: out <= 12'h222;
      20'h0798a: out <= 12'h222;
      20'h0798b: out <= 12'h222;
      20'h0798c: out <= 12'h222;
      20'h0798d: out <= 12'h222;
      20'h0798e: out <= 12'h222;
      20'h0798f: out <= 12'h222;
      20'h07990: out <= 12'h222;
      20'h07991: out <= 12'h222;
      20'h07992: out <= 12'h222;
      20'h07993: out <= 12'h222;
      20'h07994: out <= 12'h222;
      20'h07995: out <= 12'h222;
      20'h07996: out <= 12'h222;
      20'h07997: out <= 12'h222;
      20'h07998: out <= 12'h000;
      20'h07999: out <= 12'h000;
      20'h0799a: out <= 12'h000;
      20'h0799b: out <= 12'h000;
      20'h0799c: out <= 12'h000;
      20'h0799d: out <= 12'h000;
      20'h0799e: out <= 12'h000;
      20'h0799f: out <= 12'h000;
      20'h079a0: out <= 12'h000;
      20'h079a1: out <= 12'h000;
      20'h079a2: out <= 12'h000;
      20'h079a3: out <= 12'h000;
      20'h079a4: out <= 12'h000;
      20'h079a5: out <= 12'h000;
      20'h079a6: out <= 12'h000;
      20'h079a7: out <= 12'h000;
      20'h079a8: out <= 12'h222;
      20'h079a9: out <= 12'h222;
      20'h079aa: out <= 12'h222;
      20'h079ab: out <= 12'h222;
      20'h079ac: out <= 12'h222;
      20'h079ad: out <= 12'h222;
      20'h079ae: out <= 12'h222;
      20'h079af: out <= 12'h222;
      20'h079b0: out <= 12'h222;
      20'h079b1: out <= 12'h222;
      20'h079b2: out <= 12'h222;
      20'h079b3: out <= 12'h222;
      20'h079b4: out <= 12'h222;
      20'h079b5: out <= 12'h222;
      20'h079b6: out <= 12'h222;
      20'h079b7: out <= 12'h222;
      20'h079b8: out <= 12'h000;
      20'h079b9: out <= 12'h000;
      20'h079ba: out <= 12'h000;
      20'h079bb: out <= 12'h000;
      20'h079bc: out <= 12'h000;
      20'h079bd: out <= 12'h000;
      20'h079be: out <= 12'h000;
      20'h079bf: out <= 12'h000;
      20'h079c0: out <= 12'h000;
      20'h079c1: out <= 12'h000;
      20'h079c2: out <= 12'h000;
      20'h079c3: out <= 12'h000;
      20'h079c4: out <= 12'h000;
      20'h079c5: out <= 12'h000;
      20'h079c6: out <= 12'h000;
      20'h079c7: out <= 12'h000;
      20'h079c8: out <= 12'h222;
      20'h079c9: out <= 12'h222;
      20'h079ca: out <= 12'h222;
      20'h079cb: out <= 12'h222;
      20'h079cc: out <= 12'h222;
      20'h079cd: out <= 12'h222;
      20'h079ce: out <= 12'h666;
      20'h079cf: out <= 12'hbbb;
      20'h079d0: out <= 12'hfff;
      20'h079d1: out <= 12'hbbb;
      20'h079d2: out <= 12'h666;
      20'h079d3: out <= 12'h222;
      20'h079d4: out <= 12'h222;
      20'h079d5: out <= 12'h222;
      20'h079d6: out <= 12'h222;
      20'h079d7: out <= 12'h222;
      20'h079d8: out <= 12'h000;
      20'h079d9: out <= 12'h000;
      20'h079da: out <= 12'h000;
      20'h079db: out <= 12'h000;
      20'h079dc: out <= 12'h000;
      20'h079dd: out <= 12'h000;
      20'h079de: out <= 12'h666;
      20'h079df: out <= 12'hbbb;
      20'h079e0: out <= 12'hfff;
      20'h079e1: out <= 12'hbbb;
      20'h079e2: out <= 12'h666;
      20'h079e3: out <= 12'h000;
      20'h079e4: out <= 12'h000;
      20'h079e5: out <= 12'h000;
      20'h079e6: out <= 12'h000;
      20'h079e7: out <= 12'h000;
      20'h079e8: out <= 12'h603;
      20'h079e9: out <= 12'h603;
      20'h079ea: out <= 12'h603;
      20'h079eb: out <= 12'h603;
      20'h079ec: out <= 12'h603;
      20'h079ed: out <= 12'h603;
      20'h079ee: out <= 12'h603;
      20'h079ef: out <= 12'h603;
      20'h079f0: out <= 12'h603;
      20'h079f1: out <= 12'h603;
      20'h079f2: out <= 12'h603;
      20'h079f3: out <= 12'h603;
      20'h079f4: out <= 12'hb27;
      20'h079f5: out <= 12'hb27;
      20'h079f6: out <= 12'hb27;
      20'h079f7: out <= 12'hb27;
      20'h079f8: out <= 12'hb27;
      20'h079f9: out <= 12'hb27;
      20'h079fa: out <= 12'hb27;
      20'h079fb: out <= 12'hb27;
      20'h079fc: out <= 12'h603;
      20'h079fd: out <= 12'h603;
      20'h079fe: out <= 12'h603;
      20'h079ff: out <= 12'h603;
      20'h07a00: out <= 12'h603;
      20'h07a01: out <= 12'h603;
      20'h07a02: out <= 12'h603;
      20'h07a03: out <= 12'h603;
      20'h07a04: out <= 12'h603;
      20'h07a05: out <= 12'h603;
      20'h07a06: out <= 12'h603;
      20'h07a07: out <= 12'h603;
      20'h07a08: out <= 12'h603;
      20'h07a09: out <= 12'h603;
      20'h07a0a: out <= 12'h603;
      20'h07a0b: out <= 12'h603;
      20'h07a0c: out <= 12'hb27;
      20'h07a0d: out <= 12'hb27;
      20'h07a0e: out <= 12'hb27;
      20'h07a0f: out <= 12'hb27;
      20'h07a10: out <= 12'hb27;
      20'h07a11: out <= 12'hb27;
      20'h07a12: out <= 12'hb27;
      20'h07a13: out <= 12'hb27;
      20'h07a14: out <= 12'h603;
      20'h07a15: out <= 12'h603;
      20'h07a16: out <= 12'h603;
      20'h07a17: out <= 12'h603;
      20'h07a18: out <= 12'h603;
      20'h07a19: out <= 12'h603;
      20'h07a1a: out <= 12'h603;
      20'h07a1b: out <= 12'h603;
      20'h07a1c: out <= 12'h603;
      20'h07a1d: out <= 12'h603;
      20'h07a1e: out <= 12'h603;
      20'h07a1f: out <= 12'h603;
      20'h07a20: out <= 12'h603;
      20'h07a21: out <= 12'h603;
      20'h07a22: out <= 12'h603;
      20'h07a23: out <= 12'h603;
      20'h07a24: out <= 12'h603;
      20'h07a25: out <= 12'h603;
      20'h07a26: out <= 12'h603;
      20'h07a27: out <= 12'h603;
      20'h07a28: out <= 12'h603;
      20'h07a29: out <= 12'h603;
      20'h07a2a: out <= 12'h603;
      20'h07a2b: out <= 12'h603;
      20'h07a2c: out <= 12'h603;
      20'h07a2d: out <= 12'h603;
      20'h07a2e: out <= 12'h603;
      20'h07a2f: out <= 12'h603;
      20'h07a30: out <= 12'h603;
      20'h07a31: out <= 12'h603;
      20'h07a32: out <= 12'h603;
      20'h07a33: out <= 12'h603;
      20'h07a34: out <= 12'h603;
      20'h07a35: out <= 12'h603;
      20'h07a36: out <= 12'h603;
      20'h07a37: out <= 12'h603;
      20'h07a38: out <= 12'h603;
      20'h07a39: out <= 12'h603;
      20'h07a3a: out <= 12'h603;
      20'h07a3b: out <= 12'h603;
      20'h07a3c: out <= 12'h603;
      20'h07a3d: out <= 12'h603;
      20'h07a3e: out <= 12'h603;
      20'h07a3f: out <= 12'h603;
      20'h07a40: out <= 12'hb27;
      20'h07a41: out <= 12'hb27;
      20'h07a42: out <= 12'hb27;
      20'h07a43: out <= 12'hb27;
      20'h07a44: out <= 12'hb27;
      20'h07a45: out <= 12'hb27;
      20'h07a46: out <= 12'hb27;
      20'h07a47: out <= 12'hb27;
      20'h07a48: out <= 12'h000;
      20'h07a49: out <= 12'h000;
      20'h07a4a: out <= 12'h000;
      20'h07a4b: out <= 12'h000;
      20'h07a4c: out <= 12'h000;
      20'h07a4d: out <= 12'h000;
      20'h07a4e: out <= 12'h000;
      20'h07a4f: out <= 12'h000;
      20'h07a50: out <= 12'h777;
      20'h07a51: out <= 12'h777;
      20'h07a52: out <= 12'h777;
      20'h07a53: out <= 12'h777;
      20'h07a54: out <= 12'h777;
      20'h07a55: out <= 12'h777;
      20'h07a56: out <= 12'h777;
      20'h07a57: out <= 12'h777;
      20'h07a58: out <= 12'h777;
      20'h07a59: out <= 12'h777;
      20'h07a5a: out <= 12'h777;
      20'h07a5b: out <= 12'h777;
      20'h07a5c: out <= 12'h777;
      20'h07a5d: out <= 12'h777;
      20'h07a5e: out <= 12'h777;
      20'h07a5f: out <= 12'h777;
      20'h07a60: out <= 12'h000;
      20'h07a61: out <= 12'h000;
      20'h07a62: out <= 12'h000;
      20'h07a63: out <= 12'h000;
      20'h07a64: out <= 12'h000;
      20'h07a65: out <= 12'h000;
      20'h07a66: out <= 12'h000;
      20'h07a67: out <= 12'h000;
      20'h07a68: out <= 12'hfa9;
      20'h07a69: out <= 12'hfa9;
      20'h07a6a: out <= 12'hfa9;
      20'h07a6b: out <= 12'hfa9;
      20'h07a6c: out <= 12'hfa9;
      20'h07a6d: out <= 12'hfa9;
      20'h07a6e: out <= 12'hfa9;
      20'h07a6f: out <= 12'hfa9;
      20'h07a70: out <= 12'hf76;
      20'h07a71: out <= 12'hf76;
      20'h07a72: out <= 12'hf76;
      20'h07a73: out <= 12'hf76;
      20'h07a74: out <= 12'hf76;
      20'h07a75: out <= 12'hf76;
      20'h07a76: out <= 12'hf76;
      20'h07a77: out <= 12'hf76;
      20'h07a78: out <= 12'h000;
      20'h07a79: out <= 12'h000;
      20'h07a7a: out <= 12'h000;
      20'h07a7b: out <= 12'h000;
      20'h07a7c: out <= 12'h000;
      20'h07a7d: out <= 12'h000;
      20'h07a7e: out <= 12'h000;
      20'h07a7f: out <= 12'h000;
      20'h07a80: out <= 12'h000;
      20'h07a81: out <= 12'h000;
      20'h07a82: out <= 12'h000;
      20'h07a83: out <= 12'h000;
      20'h07a84: out <= 12'h000;
      20'h07a85: out <= 12'h000;
      20'h07a86: out <= 12'h000;
      20'h07a87: out <= 12'h000;
      20'h07a88: out <= 12'h000;
      20'h07a89: out <= 12'h000;
      20'h07a8a: out <= 12'h000;
      20'h07a8b: out <= 12'h000;
      20'h07a8c: out <= 12'h000;
      20'h07a8d: out <= 12'h000;
      20'h07a8e: out <= 12'h000;
      20'h07a8f: out <= 12'h000;
      20'h07a90: out <= 12'h222;
      20'h07a91: out <= 12'h222;
      20'h07a92: out <= 12'h222;
      20'h07a93: out <= 12'h222;
      20'h07a94: out <= 12'h222;
      20'h07a95: out <= 12'h222;
      20'h07a96: out <= 12'h222;
      20'h07a97: out <= 12'h222;
      20'h07a98: out <= 12'h222;
      20'h07a99: out <= 12'h222;
      20'h07a9a: out <= 12'h222;
      20'h07a9b: out <= 12'h222;
      20'h07a9c: out <= 12'h222;
      20'h07a9d: out <= 12'h222;
      20'h07a9e: out <= 12'h222;
      20'h07a9f: out <= 12'h222;
      20'h07aa0: out <= 12'h000;
      20'h07aa1: out <= 12'h000;
      20'h07aa2: out <= 12'h000;
      20'h07aa3: out <= 12'h000;
      20'h07aa4: out <= 12'h000;
      20'h07aa5: out <= 12'h000;
      20'h07aa6: out <= 12'h000;
      20'h07aa7: out <= 12'h660;
      20'h07aa8: out <= 12'hee9;
      20'h07aa9: out <= 12'h660;
      20'h07aaa: out <= 12'h000;
      20'h07aab: out <= 12'h000;
      20'h07aac: out <= 12'h000;
      20'h07aad: out <= 12'h000;
      20'h07aae: out <= 12'h000;
      20'h07aaf: out <= 12'h000;
      20'h07ab0: out <= 12'h222;
      20'h07ab1: out <= 12'h222;
      20'h07ab2: out <= 12'h222;
      20'h07ab3: out <= 12'h222;
      20'h07ab4: out <= 12'h222;
      20'h07ab5: out <= 12'h222;
      20'h07ab6: out <= 12'h222;
      20'h07ab7: out <= 12'h660;
      20'h07ab8: out <= 12'hee9;
      20'h07ab9: out <= 12'h660;
      20'h07aba: out <= 12'h222;
      20'h07abb: out <= 12'h222;
      20'h07abc: out <= 12'h222;
      20'h07abd: out <= 12'h222;
      20'h07abe: out <= 12'h222;
      20'h07abf: out <= 12'h222;
      20'h07ac0: out <= 12'h000;
      20'h07ac1: out <= 12'h000;
      20'h07ac2: out <= 12'h000;
      20'h07ac3: out <= 12'h000;
      20'h07ac4: out <= 12'h000;
      20'h07ac5: out <= 12'h000;
      20'h07ac6: out <= 12'h000;
      20'h07ac7: out <= 12'h000;
      20'h07ac8: out <= 12'h000;
      20'h07ac9: out <= 12'h000;
      20'h07aca: out <= 12'h000;
      20'h07acb: out <= 12'h000;
      20'h07acc: out <= 12'h000;
      20'h07acd: out <= 12'h000;
      20'h07ace: out <= 12'h000;
      20'h07acf: out <= 12'h000;
      20'h07ad0: out <= 12'h222;
      20'h07ad1: out <= 12'h222;
      20'h07ad2: out <= 12'h222;
      20'h07ad3: out <= 12'h222;
      20'h07ad4: out <= 12'h222;
      20'h07ad5: out <= 12'h222;
      20'h07ad6: out <= 12'h222;
      20'h07ad7: out <= 12'h222;
      20'h07ad8: out <= 12'h222;
      20'h07ad9: out <= 12'h222;
      20'h07ada: out <= 12'h222;
      20'h07adb: out <= 12'h222;
      20'h07adc: out <= 12'h222;
      20'h07add: out <= 12'h222;
      20'h07ade: out <= 12'h222;
      20'h07adf: out <= 12'h222;
      20'h07ae0: out <= 12'h000;
      20'h07ae1: out <= 12'h000;
      20'h07ae2: out <= 12'h000;
      20'h07ae3: out <= 12'h000;
      20'h07ae4: out <= 12'h000;
      20'h07ae5: out <= 12'h000;
      20'h07ae6: out <= 12'h000;
      20'h07ae7: out <= 12'h000;
      20'h07ae8: out <= 12'h000;
      20'h07ae9: out <= 12'h000;
      20'h07aea: out <= 12'h000;
      20'h07aeb: out <= 12'h000;
      20'h07aec: out <= 12'h000;
      20'h07aed: out <= 12'h000;
      20'h07aee: out <= 12'h000;
      20'h07aef: out <= 12'h000;
      20'h07af0: out <= 12'h222;
      20'h07af1: out <= 12'h222;
      20'h07af2: out <= 12'h222;
      20'h07af3: out <= 12'h222;
      20'h07af4: out <= 12'h222;
      20'h07af5: out <= 12'h222;
      20'h07af6: out <= 12'h222;
      20'h07af7: out <= 12'h222;
      20'h07af8: out <= 12'h222;
      20'h07af9: out <= 12'h222;
      20'h07afa: out <= 12'h222;
      20'h07afb: out <= 12'h222;
      20'h07afc: out <= 12'h222;
      20'h07afd: out <= 12'h222;
      20'h07afe: out <= 12'h222;
      20'h07aff: out <= 12'h222;
      20'h07b00: out <= 12'h603;
      20'h07b01: out <= 12'h603;
      20'h07b02: out <= 12'h603;
      20'h07b03: out <= 12'h603;
      20'h07b04: out <= 12'h603;
      20'h07b05: out <= 12'h603;
      20'h07b06: out <= 12'h603;
      20'h07b07: out <= 12'h603;
      20'h07b08: out <= 12'h603;
      20'h07b09: out <= 12'h603;
      20'h07b0a: out <= 12'h603;
      20'h07b0b: out <= 12'h603;
      20'h07b0c: out <= 12'hee9;
      20'h07b0d: out <= 12'hee9;
      20'h07b0e: out <= 12'hee9;
      20'h07b0f: out <= 12'hee9;
      20'h07b10: out <= 12'hee9;
      20'h07b11: out <= 12'hee9;
      20'h07b12: out <= 12'hee9;
      20'h07b13: out <= 12'hb27;
      20'h07b14: out <= 12'h603;
      20'h07b15: out <= 12'h603;
      20'h07b16: out <= 12'h603;
      20'h07b17: out <= 12'h603;
      20'h07b18: out <= 12'h603;
      20'h07b19: out <= 12'h603;
      20'h07b1a: out <= 12'h603;
      20'h07b1b: out <= 12'h603;
      20'h07b1c: out <= 12'h603;
      20'h07b1d: out <= 12'h603;
      20'h07b1e: out <= 12'h603;
      20'h07b1f: out <= 12'h603;
      20'h07b20: out <= 12'h603;
      20'h07b21: out <= 12'h603;
      20'h07b22: out <= 12'h603;
      20'h07b23: out <= 12'h603;
      20'h07b24: out <= 12'hee9;
      20'h07b25: out <= 12'hee9;
      20'h07b26: out <= 12'hee9;
      20'h07b27: out <= 12'hee9;
      20'h07b28: out <= 12'hee9;
      20'h07b29: out <= 12'hee9;
      20'h07b2a: out <= 12'hee9;
      20'h07b2b: out <= 12'hb27;
      20'h07b2c: out <= 12'h603;
      20'h07b2d: out <= 12'h603;
      20'h07b2e: out <= 12'h603;
      20'h07b2f: out <= 12'h603;
      20'h07b30: out <= 12'h603;
      20'h07b31: out <= 12'h603;
      20'h07b32: out <= 12'h603;
      20'h07b33: out <= 12'h603;
      20'h07b34: out <= 12'h603;
      20'h07b35: out <= 12'h603;
      20'h07b36: out <= 12'h603;
      20'h07b37: out <= 12'h603;
      20'h07b38: out <= 12'h603;
      20'h07b39: out <= 12'h603;
      20'h07b3a: out <= 12'h603;
      20'h07b3b: out <= 12'h603;
      20'h07b3c: out <= 12'h603;
      20'h07b3d: out <= 12'h603;
      20'h07b3e: out <= 12'h603;
      20'h07b3f: out <= 12'h603;
      20'h07b40: out <= 12'h603;
      20'h07b41: out <= 12'h603;
      20'h07b42: out <= 12'h603;
      20'h07b43: out <= 12'h603;
      20'h07b44: out <= 12'h603;
      20'h07b45: out <= 12'h603;
      20'h07b46: out <= 12'h603;
      20'h07b47: out <= 12'h603;
      20'h07b48: out <= 12'h603;
      20'h07b49: out <= 12'h603;
      20'h07b4a: out <= 12'h603;
      20'h07b4b: out <= 12'h603;
      20'h07b4c: out <= 12'h603;
      20'h07b4d: out <= 12'h603;
      20'h07b4e: out <= 12'h603;
      20'h07b4f: out <= 12'h603;
      20'h07b50: out <= 12'h603;
      20'h07b51: out <= 12'h603;
      20'h07b52: out <= 12'h603;
      20'h07b53: out <= 12'h603;
      20'h07b54: out <= 12'h603;
      20'h07b55: out <= 12'h603;
      20'h07b56: out <= 12'h603;
      20'h07b57: out <= 12'h603;
      20'h07b58: out <= 12'hee9;
      20'h07b59: out <= 12'hee9;
      20'h07b5a: out <= 12'hee9;
      20'h07b5b: out <= 12'hee9;
      20'h07b5c: out <= 12'hee9;
      20'h07b5d: out <= 12'hee9;
      20'h07b5e: out <= 12'hee9;
      20'h07b5f: out <= 12'hb27;
      20'h07b60: out <= 12'hee9;
      20'h07b61: out <= 12'hee9;
      20'h07b62: out <= 12'hee9;
      20'h07b63: out <= 12'hee9;
      20'h07b64: out <= 12'hee9;
      20'h07b65: out <= 12'hee9;
      20'h07b66: out <= 12'hee9;
      20'h07b67: out <= 12'hb27;
      20'h07b68: out <= 12'hee9;
      20'h07b69: out <= 12'hee9;
      20'h07b6a: out <= 12'hee9;
      20'h07b6b: out <= 12'hee9;
      20'h07b6c: out <= 12'hee9;
      20'h07b6d: out <= 12'hee9;
      20'h07b6e: out <= 12'hee9;
      20'h07b6f: out <= 12'hb27;
      20'h07b70: out <= 12'hee9;
      20'h07b71: out <= 12'hee9;
      20'h07b72: out <= 12'hee9;
      20'h07b73: out <= 12'hee9;
      20'h07b74: out <= 12'hee9;
      20'h07b75: out <= 12'hee9;
      20'h07b76: out <= 12'hee9;
      20'h07b77: out <= 12'hb27;
      20'h07b78: out <= 12'hee9;
      20'h07b79: out <= 12'hee9;
      20'h07b7a: out <= 12'hee9;
      20'h07b7b: out <= 12'hee9;
      20'h07b7c: out <= 12'hee9;
      20'h07b7d: out <= 12'hee9;
      20'h07b7e: out <= 12'hee9;
      20'h07b7f: out <= 12'hb27;
      20'h07b80: out <= 12'hee9;
      20'h07b81: out <= 12'hee9;
      20'h07b82: out <= 12'hee9;
      20'h07b83: out <= 12'hee9;
      20'h07b84: out <= 12'hee9;
      20'h07b85: out <= 12'hee9;
      20'h07b86: out <= 12'hee9;
      20'h07b87: out <= 12'hb27;
      20'h07b88: out <= 12'hee9;
      20'h07b89: out <= 12'hee9;
      20'h07b8a: out <= 12'hee9;
      20'h07b8b: out <= 12'hee9;
      20'h07b8c: out <= 12'hee9;
      20'h07b8d: out <= 12'hee9;
      20'h07b8e: out <= 12'hee9;
      20'h07b8f: out <= 12'hb27;
      20'h07b90: out <= 12'hee9;
      20'h07b91: out <= 12'hee9;
      20'h07b92: out <= 12'hee9;
      20'h07b93: out <= 12'hee9;
      20'h07b94: out <= 12'hee9;
      20'h07b95: out <= 12'hee9;
      20'h07b96: out <= 12'hee9;
      20'h07b97: out <= 12'hb27;
      20'h07b98: out <= 12'h000;
      20'h07b99: out <= 12'h000;
      20'h07b9a: out <= 12'h660;
      20'h07b9b: out <= 12'h660;
      20'h07b9c: out <= 12'h660;
      20'h07b9d: out <= 12'h660;
      20'h07b9e: out <= 12'h660;
      20'h07b9f: out <= 12'h660;
      20'h07ba0: out <= 12'h660;
      20'h07ba1: out <= 12'h660;
      20'h07ba2: out <= 12'h660;
      20'h07ba3: out <= 12'h660;
      20'h07ba4: out <= 12'h660;
      20'h07ba5: out <= 12'h660;
      20'h07ba6: out <= 12'h000;
      20'h07ba7: out <= 12'h000;
      20'h07ba8: out <= 12'h222;
      20'h07ba9: out <= 12'h222;
      20'h07baa: out <= 12'h660;
      20'h07bab: out <= 12'h660;
      20'h07bac: out <= 12'h660;
      20'h07bad: out <= 12'h660;
      20'h07bae: out <= 12'h660;
      20'h07baf: out <= 12'h660;
      20'h07bb0: out <= 12'h660;
      20'h07bb1: out <= 12'h660;
      20'h07bb2: out <= 12'h660;
      20'h07bb3: out <= 12'h660;
      20'h07bb4: out <= 12'h660;
      20'h07bb5: out <= 12'h660;
      20'h07bb6: out <= 12'h222;
      20'h07bb7: out <= 12'h222;
      20'h07bb8: out <= 12'h000;
      20'h07bb9: out <= 12'h000;
      20'h07bba: out <= 12'h000;
      20'h07bbb: out <= 12'h000;
      20'h07bbc: out <= 12'h000;
      20'h07bbd: out <= 12'h660;
      20'h07bbe: out <= 12'hbb0;
      20'h07bbf: out <= 12'h660;
      20'h07bc0: out <= 12'hee9;
      20'h07bc1: out <= 12'h660;
      20'h07bc2: out <= 12'hbb0;
      20'h07bc3: out <= 12'h660;
      20'h07bc4: out <= 12'h000;
      20'h07bc5: out <= 12'h000;
      20'h07bc6: out <= 12'h000;
      20'h07bc7: out <= 12'h000;
      20'h07bc8: out <= 12'h222;
      20'h07bc9: out <= 12'h222;
      20'h07bca: out <= 12'h222;
      20'h07bcb: out <= 12'h222;
      20'h07bcc: out <= 12'h222;
      20'h07bcd: out <= 12'h660;
      20'h07bce: out <= 12'hbb0;
      20'h07bcf: out <= 12'h660;
      20'h07bd0: out <= 12'hee9;
      20'h07bd1: out <= 12'h660;
      20'h07bd2: out <= 12'hbb0;
      20'h07bd3: out <= 12'h660;
      20'h07bd4: out <= 12'h222;
      20'h07bd5: out <= 12'h222;
      20'h07bd6: out <= 12'h222;
      20'h07bd7: out <= 12'h222;
      20'h07bd8: out <= 12'h000;
      20'h07bd9: out <= 12'h000;
      20'h07bda: out <= 12'h660;
      20'h07bdb: out <= 12'h660;
      20'h07bdc: out <= 12'h660;
      20'h07bdd: out <= 12'h660;
      20'h07bde: out <= 12'h660;
      20'h07bdf: out <= 12'h660;
      20'h07be0: out <= 12'h660;
      20'h07be1: out <= 12'h660;
      20'h07be2: out <= 12'h660;
      20'h07be3: out <= 12'h660;
      20'h07be4: out <= 12'h660;
      20'h07be5: out <= 12'h660;
      20'h07be6: out <= 12'h000;
      20'h07be7: out <= 12'h000;
      20'h07be8: out <= 12'h222;
      20'h07be9: out <= 12'h222;
      20'h07bea: out <= 12'h660;
      20'h07beb: out <= 12'h660;
      20'h07bec: out <= 12'h660;
      20'h07bed: out <= 12'h660;
      20'h07bee: out <= 12'h660;
      20'h07bef: out <= 12'h660;
      20'h07bf0: out <= 12'h660;
      20'h07bf1: out <= 12'h660;
      20'h07bf2: out <= 12'h660;
      20'h07bf3: out <= 12'h660;
      20'h07bf4: out <= 12'h660;
      20'h07bf5: out <= 12'h660;
      20'h07bf6: out <= 12'h222;
      20'h07bf7: out <= 12'h222;
      20'h07bf8: out <= 12'h000;
      20'h07bf9: out <= 12'h000;
      20'h07bfa: out <= 12'h000;
      20'h07bfb: out <= 12'h000;
      20'h07bfc: out <= 12'h000;
      20'h07bfd: out <= 12'h660;
      20'h07bfe: out <= 12'hbb0;
      20'h07bff: out <= 12'hbb0;
      20'h07c00: out <= 12'hbb0;
      20'h07c01: out <= 12'hbb0;
      20'h07c02: out <= 12'hbb0;
      20'h07c03: out <= 12'h660;
      20'h07c04: out <= 12'h000;
      20'h07c05: out <= 12'h000;
      20'h07c06: out <= 12'h000;
      20'h07c07: out <= 12'h000;
      20'h07c08: out <= 12'h222;
      20'h07c09: out <= 12'h222;
      20'h07c0a: out <= 12'h222;
      20'h07c0b: out <= 12'h222;
      20'h07c0c: out <= 12'h222;
      20'h07c0d: out <= 12'h660;
      20'h07c0e: out <= 12'hbb0;
      20'h07c0f: out <= 12'hbb0;
      20'h07c10: out <= 12'hbb0;
      20'h07c11: out <= 12'hbb0;
      20'h07c12: out <= 12'hbb0;
      20'h07c13: out <= 12'h660;
      20'h07c14: out <= 12'h222;
      20'h07c15: out <= 12'h222;
      20'h07c16: out <= 12'h222;
      20'h07c17: out <= 12'h222;
      20'h07c18: out <= 12'h603;
      20'h07c19: out <= 12'h603;
      20'h07c1a: out <= 12'h603;
      20'h07c1b: out <= 12'h603;
      20'h07c1c: out <= 12'h603;
      20'h07c1d: out <= 12'h603;
      20'h07c1e: out <= 12'h603;
      20'h07c1f: out <= 12'h603;
      20'h07c20: out <= 12'h603;
      20'h07c21: out <= 12'h603;
      20'h07c22: out <= 12'h603;
      20'h07c23: out <= 12'h603;
      20'h07c24: out <= 12'hee9;
      20'h07c25: out <= 12'hf87;
      20'h07c26: out <= 12'hf87;
      20'h07c27: out <= 12'hf87;
      20'h07c28: out <= 12'hf87;
      20'h07c29: out <= 12'hf87;
      20'h07c2a: out <= 12'hf87;
      20'h07c2b: out <= 12'hb27;
      20'h07c2c: out <= 12'h603;
      20'h07c2d: out <= 12'h603;
      20'h07c2e: out <= 12'h603;
      20'h07c2f: out <= 12'h603;
      20'h07c30: out <= 12'h603;
      20'h07c31: out <= 12'h603;
      20'h07c32: out <= 12'h603;
      20'h07c33: out <= 12'h603;
      20'h07c34: out <= 12'h603;
      20'h07c35: out <= 12'h603;
      20'h07c36: out <= 12'h603;
      20'h07c37: out <= 12'h603;
      20'h07c38: out <= 12'h603;
      20'h07c39: out <= 12'h603;
      20'h07c3a: out <= 12'h603;
      20'h07c3b: out <= 12'h603;
      20'h07c3c: out <= 12'hee9;
      20'h07c3d: out <= 12'hf87;
      20'h07c3e: out <= 12'hf87;
      20'h07c3f: out <= 12'hf87;
      20'h07c40: out <= 12'hf87;
      20'h07c41: out <= 12'hf87;
      20'h07c42: out <= 12'hf87;
      20'h07c43: out <= 12'hb27;
      20'h07c44: out <= 12'h603;
      20'h07c45: out <= 12'h603;
      20'h07c46: out <= 12'h603;
      20'h07c47: out <= 12'h603;
      20'h07c48: out <= 12'h603;
      20'h07c49: out <= 12'h603;
      20'h07c4a: out <= 12'h603;
      20'h07c4b: out <= 12'h603;
      20'h07c4c: out <= 12'h603;
      20'h07c4d: out <= 12'h603;
      20'h07c4e: out <= 12'h603;
      20'h07c4f: out <= 12'h603;
      20'h07c50: out <= 12'h603;
      20'h07c51: out <= 12'h603;
      20'h07c52: out <= 12'h603;
      20'h07c53: out <= 12'h603;
      20'h07c54: out <= 12'h603;
      20'h07c55: out <= 12'h603;
      20'h07c56: out <= 12'h603;
      20'h07c57: out <= 12'h603;
      20'h07c58: out <= 12'h603;
      20'h07c59: out <= 12'h603;
      20'h07c5a: out <= 12'h603;
      20'h07c5b: out <= 12'h603;
      20'h07c5c: out <= 12'h603;
      20'h07c5d: out <= 12'h603;
      20'h07c5e: out <= 12'h603;
      20'h07c5f: out <= 12'h603;
      20'h07c60: out <= 12'h603;
      20'h07c61: out <= 12'h603;
      20'h07c62: out <= 12'h603;
      20'h07c63: out <= 12'h603;
      20'h07c64: out <= 12'h603;
      20'h07c65: out <= 12'h603;
      20'h07c66: out <= 12'h603;
      20'h07c67: out <= 12'h603;
      20'h07c68: out <= 12'h603;
      20'h07c69: out <= 12'h603;
      20'h07c6a: out <= 12'h603;
      20'h07c6b: out <= 12'h603;
      20'h07c6c: out <= 12'h603;
      20'h07c6d: out <= 12'h603;
      20'h07c6e: out <= 12'h603;
      20'h07c6f: out <= 12'h603;
      20'h07c70: out <= 12'hee9;
      20'h07c71: out <= 12'hf87;
      20'h07c72: out <= 12'hf87;
      20'h07c73: out <= 12'hf87;
      20'h07c74: out <= 12'hf87;
      20'h07c75: out <= 12'hf87;
      20'h07c76: out <= 12'hf87;
      20'h07c77: out <= 12'hb27;
      20'h07c78: out <= 12'hee9;
      20'h07c79: out <= 12'hf87;
      20'h07c7a: out <= 12'hf87;
      20'h07c7b: out <= 12'hf87;
      20'h07c7c: out <= 12'hf87;
      20'h07c7d: out <= 12'hf87;
      20'h07c7e: out <= 12'hf87;
      20'h07c7f: out <= 12'hb27;
      20'h07c80: out <= 12'hee9;
      20'h07c81: out <= 12'hf87;
      20'h07c82: out <= 12'hf87;
      20'h07c83: out <= 12'hf87;
      20'h07c84: out <= 12'hf87;
      20'h07c85: out <= 12'hf87;
      20'h07c86: out <= 12'hf87;
      20'h07c87: out <= 12'hb27;
      20'h07c88: out <= 12'hee9;
      20'h07c89: out <= 12'hf87;
      20'h07c8a: out <= 12'hf87;
      20'h07c8b: out <= 12'hf87;
      20'h07c8c: out <= 12'hf87;
      20'h07c8d: out <= 12'hf87;
      20'h07c8e: out <= 12'hf87;
      20'h07c8f: out <= 12'hb27;
      20'h07c90: out <= 12'hee9;
      20'h07c91: out <= 12'hf87;
      20'h07c92: out <= 12'hf87;
      20'h07c93: out <= 12'hf87;
      20'h07c94: out <= 12'hf87;
      20'h07c95: out <= 12'hf87;
      20'h07c96: out <= 12'hf87;
      20'h07c97: out <= 12'hb27;
      20'h07c98: out <= 12'hee9;
      20'h07c99: out <= 12'hf87;
      20'h07c9a: out <= 12'hf87;
      20'h07c9b: out <= 12'hf87;
      20'h07c9c: out <= 12'hf87;
      20'h07c9d: out <= 12'hf87;
      20'h07c9e: out <= 12'hf87;
      20'h07c9f: out <= 12'hb27;
      20'h07ca0: out <= 12'hee9;
      20'h07ca1: out <= 12'hf87;
      20'h07ca2: out <= 12'hf87;
      20'h07ca3: out <= 12'hf87;
      20'h07ca4: out <= 12'hf87;
      20'h07ca5: out <= 12'hf87;
      20'h07ca6: out <= 12'hf87;
      20'h07ca7: out <= 12'hb27;
      20'h07ca8: out <= 12'hee9;
      20'h07ca9: out <= 12'hf87;
      20'h07caa: out <= 12'hf87;
      20'h07cab: out <= 12'hf87;
      20'h07cac: out <= 12'hf87;
      20'h07cad: out <= 12'hf87;
      20'h07cae: out <= 12'hf87;
      20'h07caf: out <= 12'hb27;
      20'h07cb0: out <= 12'h000;
      20'h07cb1: out <= 12'h000;
      20'h07cb2: out <= 12'hee9;
      20'h07cb3: out <= 12'h660;
      20'h07cb4: out <= 12'hee9;
      20'h07cb5: out <= 12'h660;
      20'h07cb6: out <= 12'hee9;
      20'h07cb7: out <= 12'h660;
      20'h07cb8: out <= 12'hee9;
      20'h07cb9: out <= 12'h660;
      20'h07cba: out <= 12'hee9;
      20'h07cbb: out <= 12'h660;
      20'h07cbc: out <= 12'hee9;
      20'h07cbd: out <= 12'h660;
      20'h07cbe: out <= 12'h000;
      20'h07cbf: out <= 12'h000;
      20'h07cc0: out <= 12'h222;
      20'h07cc1: out <= 12'h222;
      20'h07cc2: out <= 12'h660;
      20'h07cc3: out <= 12'hee9;
      20'h07cc4: out <= 12'h660;
      20'h07cc5: out <= 12'hee9;
      20'h07cc6: out <= 12'h660;
      20'h07cc7: out <= 12'hee9;
      20'h07cc8: out <= 12'h660;
      20'h07cc9: out <= 12'hee9;
      20'h07cca: out <= 12'h660;
      20'h07ccb: out <= 12'hee9;
      20'h07ccc: out <= 12'h660;
      20'h07ccd: out <= 12'hee9;
      20'h07cce: out <= 12'h222;
      20'h07ccf: out <= 12'h222;
      20'h07cd0: out <= 12'h000;
      20'h07cd1: out <= 12'h000;
      20'h07cd2: out <= 12'h660;
      20'h07cd3: out <= 12'h660;
      20'h07cd4: out <= 12'h660;
      20'h07cd5: out <= 12'hbb0;
      20'h07cd6: out <= 12'hee9;
      20'h07cd7: out <= 12'h660;
      20'h07cd8: out <= 12'hee9;
      20'h07cd9: out <= 12'h660;
      20'h07cda: out <= 12'hee9;
      20'h07cdb: out <= 12'hbb0;
      20'h07cdc: out <= 12'h660;
      20'h07cdd: out <= 12'h660;
      20'h07cde: out <= 12'h660;
      20'h07cdf: out <= 12'h000;
      20'h07ce0: out <= 12'h222;
      20'h07ce1: out <= 12'h222;
      20'h07ce2: out <= 12'h660;
      20'h07ce3: out <= 12'hee9;
      20'h07ce4: out <= 12'h660;
      20'h07ce5: out <= 12'hbb0;
      20'h07ce6: out <= 12'hee9;
      20'h07ce7: out <= 12'h660;
      20'h07ce8: out <= 12'hee9;
      20'h07ce9: out <= 12'h660;
      20'h07cea: out <= 12'hee9;
      20'h07ceb: out <= 12'hbb0;
      20'h07cec: out <= 12'h660;
      20'h07ced: out <= 12'hee9;
      20'h07cee: out <= 12'h660;
      20'h07cef: out <= 12'h222;
      20'h07cf0: out <= 12'h000;
      20'h07cf1: out <= 12'h000;
      20'h07cf2: out <= 12'h660;
      20'h07cf3: out <= 12'hee9;
      20'h07cf4: out <= 12'h660;
      20'h07cf5: out <= 12'hee9;
      20'h07cf6: out <= 12'h660;
      20'h07cf7: out <= 12'hee9;
      20'h07cf8: out <= 12'h660;
      20'h07cf9: out <= 12'hee9;
      20'h07cfa: out <= 12'h660;
      20'h07cfb: out <= 12'hee9;
      20'h07cfc: out <= 12'h660;
      20'h07cfd: out <= 12'hee9;
      20'h07cfe: out <= 12'h000;
      20'h07cff: out <= 12'h000;
      20'h07d00: out <= 12'h222;
      20'h07d01: out <= 12'h222;
      20'h07d02: out <= 12'hee9;
      20'h07d03: out <= 12'h660;
      20'h07d04: out <= 12'hee9;
      20'h07d05: out <= 12'h660;
      20'h07d06: out <= 12'hee9;
      20'h07d07: out <= 12'h660;
      20'h07d08: out <= 12'hee9;
      20'h07d09: out <= 12'h660;
      20'h07d0a: out <= 12'hee9;
      20'h07d0b: out <= 12'h660;
      20'h07d0c: out <= 12'hee9;
      20'h07d0d: out <= 12'h660;
      20'h07d0e: out <= 12'h222;
      20'h07d0f: out <= 12'h222;
      20'h07d10: out <= 12'h000;
      20'h07d11: out <= 12'h000;
      20'h07d12: out <= 12'h660;
      20'h07d13: out <= 12'hee9;
      20'h07d14: out <= 12'h660;
      20'h07d15: out <= 12'hbb0;
      20'h07d16: out <= 12'hee9;
      20'h07d17: out <= 12'hee9;
      20'h07d18: out <= 12'hee9;
      20'h07d19: out <= 12'hee9;
      20'h07d1a: out <= 12'hee9;
      20'h07d1b: out <= 12'hbb0;
      20'h07d1c: out <= 12'h660;
      20'h07d1d: out <= 12'hee9;
      20'h07d1e: out <= 12'h660;
      20'h07d1f: out <= 12'h000;
      20'h07d20: out <= 12'h222;
      20'h07d21: out <= 12'h222;
      20'h07d22: out <= 12'h660;
      20'h07d23: out <= 12'h660;
      20'h07d24: out <= 12'h660;
      20'h07d25: out <= 12'hbb0;
      20'h07d26: out <= 12'hee9;
      20'h07d27: out <= 12'hee9;
      20'h07d28: out <= 12'hee9;
      20'h07d29: out <= 12'hee9;
      20'h07d2a: out <= 12'hee9;
      20'h07d2b: out <= 12'hbb0;
      20'h07d2c: out <= 12'h660;
      20'h07d2d: out <= 12'h660;
      20'h07d2e: out <= 12'h660;
      20'h07d2f: out <= 12'h222;
      20'h07d30: out <= 12'h603;
      20'h07d31: out <= 12'h603;
      20'h07d32: out <= 12'h603;
      20'h07d33: out <= 12'h603;
      20'h07d34: out <= 12'h603;
      20'h07d35: out <= 12'h603;
      20'h07d36: out <= 12'h603;
      20'h07d37: out <= 12'h603;
      20'h07d38: out <= 12'h603;
      20'h07d39: out <= 12'h603;
      20'h07d3a: out <= 12'h603;
      20'h07d3b: out <= 12'h603;
      20'h07d3c: out <= 12'hee9;
      20'h07d3d: out <= 12'hf87;
      20'h07d3e: out <= 12'hee9;
      20'h07d3f: out <= 12'hee9;
      20'h07d40: out <= 12'hee9;
      20'h07d41: out <= 12'hb27;
      20'h07d42: out <= 12'hf87;
      20'h07d43: out <= 12'hb27;
      20'h07d44: out <= 12'h603;
      20'h07d45: out <= 12'h603;
      20'h07d46: out <= 12'h603;
      20'h07d47: out <= 12'h603;
      20'h07d48: out <= 12'h603;
      20'h07d49: out <= 12'h603;
      20'h07d4a: out <= 12'h603;
      20'h07d4b: out <= 12'h603;
      20'h07d4c: out <= 12'h603;
      20'h07d4d: out <= 12'h603;
      20'h07d4e: out <= 12'h603;
      20'h07d4f: out <= 12'h603;
      20'h07d50: out <= 12'h603;
      20'h07d51: out <= 12'h603;
      20'h07d52: out <= 12'h603;
      20'h07d53: out <= 12'h603;
      20'h07d54: out <= 12'hee9;
      20'h07d55: out <= 12'hf87;
      20'h07d56: out <= 12'hee9;
      20'h07d57: out <= 12'hee9;
      20'h07d58: out <= 12'hee9;
      20'h07d59: out <= 12'hb27;
      20'h07d5a: out <= 12'hf87;
      20'h07d5b: out <= 12'hb27;
      20'h07d5c: out <= 12'h603;
      20'h07d5d: out <= 12'h603;
      20'h07d5e: out <= 12'h603;
      20'h07d5f: out <= 12'h603;
      20'h07d60: out <= 12'h603;
      20'h07d61: out <= 12'h603;
      20'h07d62: out <= 12'h603;
      20'h07d63: out <= 12'h603;
      20'h07d64: out <= 12'h603;
      20'h07d65: out <= 12'h603;
      20'h07d66: out <= 12'h603;
      20'h07d67: out <= 12'h603;
      20'h07d68: out <= 12'h603;
      20'h07d69: out <= 12'h603;
      20'h07d6a: out <= 12'h603;
      20'h07d6b: out <= 12'h603;
      20'h07d6c: out <= 12'h603;
      20'h07d6d: out <= 12'h603;
      20'h07d6e: out <= 12'h603;
      20'h07d6f: out <= 12'h603;
      20'h07d70: out <= 12'h603;
      20'h07d71: out <= 12'h603;
      20'h07d72: out <= 12'h603;
      20'h07d73: out <= 12'h603;
      20'h07d74: out <= 12'h603;
      20'h07d75: out <= 12'h603;
      20'h07d76: out <= 12'h603;
      20'h07d77: out <= 12'h603;
      20'h07d78: out <= 12'h603;
      20'h07d79: out <= 12'h603;
      20'h07d7a: out <= 12'h603;
      20'h07d7b: out <= 12'h603;
      20'h07d7c: out <= 12'h603;
      20'h07d7d: out <= 12'h603;
      20'h07d7e: out <= 12'h603;
      20'h07d7f: out <= 12'h603;
      20'h07d80: out <= 12'h603;
      20'h07d81: out <= 12'h603;
      20'h07d82: out <= 12'h603;
      20'h07d83: out <= 12'h603;
      20'h07d84: out <= 12'h603;
      20'h07d85: out <= 12'h603;
      20'h07d86: out <= 12'h603;
      20'h07d87: out <= 12'h603;
      20'h07d88: out <= 12'hee9;
      20'h07d89: out <= 12'hf87;
      20'h07d8a: out <= 12'hee9;
      20'h07d8b: out <= 12'hee9;
      20'h07d8c: out <= 12'hee9;
      20'h07d8d: out <= 12'hb27;
      20'h07d8e: out <= 12'hf87;
      20'h07d8f: out <= 12'hb27;
      20'h07d90: out <= 12'hee9;
      20'h07d91: out <= 12'hf87;
      20'h07d92: out <= 12'hee9;
      20'h07d93: out <= 12'hee9;
      20'h07d94: out <= 12'hee9;
      20'h07d95: out <= 12'hb27;
      20'h07d96: out <= 12'hf87;
      20'h07d97: out <= 12'hb27;
      20'h07d98: out <= 12'hee9;
      20'h07d99: out <= 12'hf87;
      20'h07d9a: out <= 12'hee9;
      20'h07d9b: out <= 12'hee9;
      20'h07d9c: out <= 12'hee9;
      20'h07d9d: out <= 12'hb27;
      20'h07d9e: out <= 12'hf87;
      20'h07d9f: out <= 12'hb27;
      20'h07da0: out <= 12'hee9;
      20'h07da1: out <= 12'hf87;
      20'h07da2: out <= 12'hee9;
      20'h07da3: out <= 12'hee9;
      20'h07da4: out <= 12'hee9;
      20'h07da5: out <= 12'hb27;
      20'h07da6: out <= 12'hf87;
      20'h07da7: out <= 12'hb27;
      20'h07da8: out <= 12'hee9;
      20'h07da9: out <= 12'hf87;
      20'h07daa: out <= 12'hee9;
      20'h07dab: out <= 12'hee9;
      20'h07dac: out <= 12'hee9;
      20'h07dad: out <= 12'hb27;
      20'h07dae: out <= 12'hf87;
      20'h07daf: out <= 12'hb27;
      20'h07db0: out <= 12'hee9;
      20'h07db1: out <= 12'hf87;
      20'h07db2: out <= 12'hee9;
      20'h07db3: out <= 12'hee9;
      20'h07db4: out <= 12'hee9;
      20'h07db5: out <= 12'hb27;
      20'h07db6: out <= 12'hf87;
      20'h07db7: out <= 12'hb27;
      20'h07db8: out <= 12'hee9;
      20'h07db9: out <= 12'hf87;
      20'h07dba: out <= 12'hee9;
      20'h07dbb: out <= 12'hee9;
      20'h07dbc: out <= 12'hee9;
      20'h07dbd: out <= 12'hb27;
      20'h07dbe: out <= 12'hf87;
      20'h07dbf: out <= 12'hb27;
      20'h07dc0: out <= 12'hee9;
      20'h07dc1: out <= 12'hf87;
      20'h07dc2: out <= 12'hee9;
      20'h07dc3: out <= 12'hee9;
      20'h07dc4: out <= 12'hee9;
      20'h07dc5: out <= 12'hb27;
      20'h07dc6: out <= 12'hf87;
      20'h07dc7: out <= 12'hb27;
      20'h07dc8: out <= 12'h000;
      20'h07dc9: out <= 12'h000;
      20'h07dca: out <= 12'h660;
      20'h07dcb: out <= 12'hbb0;
      20'h07dcc: out <= 12'hbb0;
      20'h07dcd: out <= 12'hbb0;
      20'h07dce: out <= 12'hbb0;
      20'h07dcf: out <= 12'hbb0;
      20'h07dd0: out <= 12'hbb0;
      20'h07dd1: out <= 12'hbb0;
      20'h07dd2: out <= 12'hbb0;
      20'h07dd3: out <= 12'hbb0;
      20'h07dd4: out <= 12'hbb0;
      20'h07dd5: out <= 12'h660;
      20'h07dd6: out <= 12'h000;
      20'h07dd7: out <= 12'h000;
      20'h07dd8: out <= 12'h222;
      20'h07dd9: out <= 12'h222;
      20'h07dda: out <= 12'h660;
      20'h07ddb: out <= 12'hbb0;
      20'h07ddc: out <= 12'hbb0;
      20'h07ddd: out <= 12'hbb0;
      20'h07dde: out <= 12'hbb0;
      20'h07ddf: out <= 12'hbb0;
      20'h07de0: out <= 12'hbb0;
      20'h07de1: out <= 12'hbb0;
      20'h07de2: out <= 12'hbb0;
      20'h07de3: out <= 12'hbb0;
      20'h07de4: out <= 12'hbb0;
      20'h07de5: out <= 12'h660;
      20'h07de6: out <= 12'h222;
      20'h07de7: out <= 12'h222;
      20'h07de8: out <= 12'h000;
      20'h07de9: out <= 12'h000;
      20'h07dea: out <= 12'h660;
      20'h07deb: out <= 12'hee9;
      20'h07dec: out <= 12'hbb0;
      20'h07ded: out <= 12'hee9;
      20'h07dee: out <= 12'h660;
      20'h07def: out <= 12'h660;
      20'h07df0: out <= 12'hee9;
      20'h07df1: out <= 12'h660;
      20'h07df2: out <= 12'h660;
      20'h07df3: out <= 12'hee9;
      20'h07df4: out <= 12'hbb0;
      20'h07df5: out <= 12'hee9;
      20'h07df6: out <= 12'h660;
      20'h07df7: out <= 12'h000;
      20'h07df8: out <= 12'h222;
      20'h07df9: out <= 12'h222;
      20'h07dfa: out <= 12'h660;
      20'h07dfb: out <= 12'h660;
      20'h07dfc: out <= 12'hbb0;
      20'h07dfd: out <= 12'hee9;
      20'h07dfe: out <= 12'h660;
      20'h07dff: out <= 12'h660;
      20'h07e00: out <= 12'hee9;
      20'h07e01: out <= 12'h660;
      20'h07e02: out <= 12'h660;
      20'h07e03: out <= 12'hee9;
      20'h07e04: out <= 12'hbb0;
      20'h07e05: out <= 12'h660;
      20'h07e06: out <= 12'h660;
      20'h07e07: out <= 12'h222;
      20'h07e08: out <= 12'h000;
      20'h07e09: out <= 12'h000;
      20'h07e0a: out <= 12'h660;
      20'h07e0b: out <= 12'hbb0;
      20'h07e0c: out <= 12'hbb0;
      20'h07e0d: out <= 12'hbb0;
      20'h07e0e: out <= 12'hbb0;
      20'h07e0f: out <= 12'hbb0;
      20'h07e10: out <= 12'hbb0;
      20'h07e11: out <= 12'hbb0;
      20'h07e12: out <= 12'hbb0;
      20'h07e13: out <= 12'hbb0;
      20'h07e14: out <= 12'hbb0;
      20'h07e15: out <= 12'h660;
      20'h07e16: out <= 12'h000;
      20'h07e17: out <= 12'h000;
      20'h07e18: out <= 12'h222;
      20'h07e19: out <= 12'h222;
      20'h07e1a: out <= 12'h660;
      20'h07e1b: out <= 12'hbb0;
      20'h07e1c: out <= 12'hbb0;
      20'h07e1d: out <= 12'hbb0;
      20'h07e1e: out <= 12'hbb0;
      20'h07e1f: out <= 12'hbb0;
      20'h07e20: out <= 12'hbb0;
      20'h07e21: out <= 12'hbb0;
      20'h07e22: out <= 12'hbb0;
      20'h07e23: out <= 12'hbb0;
      20'h07e24: out <= 12'hbb0;
      20'h07e25: out <= 12'h660;
      20'h07e26: out <= 12'h222;
      20'h07e27: out <= 12'h222;
      20'h07e28: out <= 12'h000;
      20'h07e29: out <= 12'h000;
      20'h07e2a: out <= 12'h660;
      20'h07e2b: out <= 12'h660;
      20'h07e2c: out <= 12'hbb0;
      20'h07e2d: out <= 12'hee9;
      20'h07e2e: out <= 12'hbb0;
      20'h07e2f: out <= 12'hbb0;
      20'h07e30: out <= 12'hbb0;
      20'h07e31: out <= 12'hbb0;
      20'h07e32: out <= 12'hbb0;
      20'h07e33: out <= 12'hee9;
      20'h07e34: out <= 12'hbb0;
      20'h07e35: out <= 12'h660;
      20'h07e36: out <= 12'h660;
      20'h07e37: out <= 12'h000;
      20'h07e38: out <= 12'h222;
      20'h07e39: out <= 12'h222;
      20'h07e3a: out <= 12'h660;
      20'h07e3b: out <= 12'hee9;
      20'h07e3c: out <= 12'hbb0;
      20'h07e3d: out <= 12'hee9;
      20'h07e3e: out <= 12'hbb0;
      20'h07e3f: out <= 12'hbb0;
      20'h07e40: out <= 12'hbb0;
      20'h07e41: out <= 12'hbb0;
      20'h07e42: out <= 12'hbb0;
      20'h07e43: out <= 12'hee9;
      20'h07e44: out <= 12'hbb0;
      20'h07e45: out <= 12'hee9;
      20'h07e46: out <= 12'h660;
      20'h07e47: out <= 12'h222;
      20'h07e48: out <= 12'h603;
      20'h07e49: out <= 12'h603;
      20'h07e4a: out <= 12'h603;
      20'h07e4b: out <= 12'h603;
      20'h07e4c: out <= 12'h603;
      20'h07e4d: out <= 12'h603;
      20'h07e4e: out <= 12'h603;
      20'h07e4f: out <= 12'h603;
      20'h07e50: out <= 12'h603;
      20'h07e51: out <= 12'h603;
      20'h07e52: out <= 12'h603;
      20'h07e53: out <= 12'h603;
      20'h07e54: out <= 12'hee9;
      20'h07e55: out <= 12'hf87;
      20'h07e56: out <= 12'hee9;
      20'h07e57: out <= 12'hf87;
      20'h07e58: out <= 12'hf87;
      20'h07e59: out <= 12'hb27;
      20'h07e5a: out <= 12'hf87;
      20'h07e5b: out <= 12'hb27;
      20'h07e5c: out <= 12'h603;
      20'h07e5d: out <= 12'h603;
      20'h07e5e: out <= 12'h603;
      20'h07e5f: out <= 12'h603;
      20'h07e60: out <= 12'h603;
      20'h07e61: out <= 12'h603;
      20'h07e62: out <= 12'h603;
      20'h07e63: out <= 12'h603;
      20'h07e64: out <= 12'h603;
      20'h07e65: out <= 12'h603;
      20'h07e66: out <= 12'h603;
      20'h07e67: out <= 12'h603;
      20'h07e68: out <= 12'h603;
      20'h07e69: out <= 12'h603;
      20'h07e6a: out <= 12'h603;
      20'h07e6b: out <= 12'h603;
      20'h07e6c: out <= 12'hee9;
      20'h07e6d: out <= 12'hf87;
      20'h07e6e: out <= 12'hee9;
      20'h07e6f: out <= 12'hf87;
      20'h07e70: out <= 12'hf87;
      20'h07e71: out <= 12'hb27;
      20'h07e72: out <= 12'hf87;
      20'h07e73: out <= 12'hb27;
      20'h07e74: out <= 12'h603;
      20'h07e75: out <= 12'h603;
      20'h07e76: out <= 12'h603;
      20'h07e77: out <= 12'h603;
      20'h07e78: out <= 12'h603;
      20'h07e79: out <= 12'h603;
      20'h07e7a: out <= 12'h603;
      20'h07e7b: out <= 12'h603;
      20'h07e7c: out <= 12'h603;
      20'h07e7d: out <= 12'h603;
      20'h07e7e: out <= 12'h603;
      20'h07e7f: out <= 12'h603;
      20'h07e80: out <= 12'h603;
      20'h07e81: out <= 12'h603;
      20'h07e82: out <= 12'h603;
      20'h07e83: out <= 12'h603;
      20'h07e84: out <= 12'h603;
      20'h07e85: out <= 12'h603;
      20'h07e86: out <= 12'h603;
      20'h07e87: out <= 12'h603;
      20'h07e88: out <= 12'h603;
      20'h07e89: out <= 12'h603;
      20'h07e8a: out <= 12'h603;
      20'h07e8b: out <= 12'h603;
      20'h07e8c: out <= 12'h603;
      20'h07e8d: out <= 12'h603;
      20'h07e8e: out <= 12'h603;
      20'h07e8f: out <= 12'h603;
      20'h07e90: out <= 12'h603;
      20'h07e91: out <= 12'h603;
      20'h07e92: out <= 12'h603;
      20'h07e93: out <= 12'h603;
      20'h07e94: out <= 12'h603;
      20'h07e95: out <= 12'h603;
      20'h07e96: out <= 12'h603;
      20'h07e97: out <= 12'h603;
      20'h07e98: out <= 12'h603;
      20'h07e99: out <= 12'h603;
      20'h07e9a: out <= 12'h603;
      20'h07e9b: out <= 12'h603;
      20'h07e9c: out <= 12'h603;
      20'h07e9d: out <= 12'h603;
      20'h07e9e: out <= 12'h603;
      20'h07e9f: out <= 12'h603;
      20'h07ea0: out <= 12'hee9;
      20'h07ea1: out <= 12'hf87;
      20'h07ea2: out <= 12'hee9;
      20'h07ea3: out <= 12'hf87;
      20'h07ea4: out <= 12'hf87;
      20'h07ea5: out <= 12'hb27;
      20'h07ea6: out <= 12'hf87;
      20'h07ea7: out <= 12'hb27;
      20'h07ea8: out <= 12'hee9;
      20'h07ea9: out <= 12'hf87;
      20'h07eaa: out <= 12'hee9;
      20'h07eab: out <= 12'hf87;
      20'h07eac: out <= 12'hf87;
      20'h07ead: out <= 12'hb27;
      20'h07eae: out <= 12'hf87;
      20'h07eaf: out <= 12'hb27;
      20'h07eb0: out <= 12'hee9;
      20'h07eb1: out <= 12'hf87;
      20'h07eb2: out <= 12'hee9;
      20'h07eb3: out <= 12'hf87;
      20'h07eb4: out <= 12'hf87;
      20'h07eb5: out <= 12'hb27;
      20'h07eb6: out <= 12'hf87;
      20'h07eb7: out <= 12'hb27;
      20'h07eb8: out <= 12'hee9;
      20'h07eb9: out <= 12'hf87;
      20'h07eba: out <= 12'hee9;
      20'h07ebb: out <= 12'hf87;
      20'h07ebc: out <= 12'hf87;
      20'h07ebd: out <= 12'hb27;
      20'h07ebe: out <= 12'hf87;
      20'h07ebf: out <= 12'hb27;
      20'h07ec0: out <= 12'hee9;
      20'h07ec1: out <= 12'hf87;
      20'h07ec2: out <= 12'hee9;
      20'h07ec3: out <= 12'hf87;
      20'h07ec4: out <= 12'hf87;
      20'h07ec5: out <= 12'hb27;
      20'h07ec6: out <= 12'hf87;
      20'h07ec7: out <= 12'hb27;
      20'h07ec8: out <= 12'hee9;
      20'h07ec9: out <= 12'hf87;
      20'h07eca: out <= 12'hee9;
      20'h07ecb: out <= 12'hf87;
      20'h07ecc: out <= 12'hf87;
      20'h07ecd: out <= 12'hb27;
      20'h07ece: out <= 12'hf87;
      20'h07ecf: out <= 12'hb27;
      20'h07ed0: out <= 12'hee9;
      20'h07ed1: out <= 12'hf87;
      20'h07ed2: out <= 12'hee9;
      20'h07ed3: out <= 12'hf87;
      20'h07ed4: out <= 12'hf87;
      20'h07ed5: out <= 12'hb27;
      20'h07ed6: out <= 12'hf87;
      20'h07ed7: out <= 12'hb27;
      20'h07ed8: out <= 12'hee9;
      20'h07ed9: out <= 12'hf87;
      20'h07eda: out <= 12'hee9;
      20'h07edb: out <= 12'hf87;
      20'h07edc: out <= 12'hf87;
      20'h07edd: out <= 12'hb27;
      20'h07ede: out <= 12'hf87;
      20'h07edf: out <= 12'hb27;
      20'h07ee0: out <= 12'h000;
      20'h07ee1: out <= 12'h660;
      20'h07ee2: out <= 12'hbb0;
      20'h07ee3: out <= 12'hee9;
      20'h07ee4: out <= 12'h660;
      20'h07ee5: out <= 12'h660;
      20'h07ee6: out <= 12'h660;
      20'h07ee7: out <= 12'h660;
      20'h07ee8: out <= 12'h660;
      20'h07ee9: out <= 12'h660;
      20'h07eea: out <= 12'hbb0;
      20'h07eeb: out <= 12'hbb0;
      20'h07eec: out <= 12'hee9;
      20'h07eed: out <= 12'hbb0;
      20'h07eee: out <= 12'h660;
      20'h07eef: out <= 12'h000;
      20'h07ef0: out <= 12'h222;
      20'h07ef1: out <= 12'h660;
      20'h07ef2: out <= 12'hbb0;
      20'h07ef3: out <= 12'hee9;
      20'h07ef4: out <= 12'h660;
      20'h07ef5: out <= 12'h660;
      20'h07ef6: out <= 12'h660;
      20'h07ef7: out <= 12'h660;
      20'h07ef8: out <= 12'h660;
      20'h07ef9: out <= 12'h660;
      20'h07efa: out <= 12'h660;
      20'h07efb: out <= 12'hbb0;
      20'h07efc: out <= 12'hee9;
      20'h07efd: out <= 12'hbb0;
      20'h07efe: out <= 12'h660;
      20'h07eff: out <= 12'h222;
      20'h07f00: out <= 12'h000;
      20'h07f01: out <= 12'h000;
      20'h07f02: out <= 12'h660;
      20'h07f03: out <= 12'h660;
      20'h07f04: out <= 12'hbb0;
      20'h07f05: out <= 12'hbb0;
      20'h07f06: out <= 12'h660;
      20'h07f07: out <= 12'hbb0;
      20'h07f08: out <= 12'hee9;
      20'h07f09: out <= 12'hbb0;
      20'h07f0a: out <= 12'h660;
      20'h07f0b: out <= 12'hbb0;
      20'h07f0c: out <= 12'hbb0;
      20'h07f0d: out <= 12'h660;
      20'h07f0e: out <= 12'h660;
      20'h07f0f: out <= 12'h000;
      20'h07f10: out <= 12'h222;
      20'h07f11: out <= 12'h222;
      20'h07f12: out <= 12'h660;
      20'h07f13: out <= 12'hee9;
      20'h07f14: out <= 12'hbb0;
      20'h07f15: out <= 12'hbb0;
      20'h07f16: out <= 12'h660;
      20'h07f17: out <= 12'hbb0;
      20'h07f18: out <= 12'hee9;
      20'h07f19: out <= 12'hbb0;
      20'h07f1a: out <= 12'h660;
      20'h07f1b: out <= 12'hbb0;
      20'h07f1c: out <= 12'hbb0;
      20'h07f1d: out <= 12'hee9;
      20'h07f1e: out <= 12'h660;
      20'h07f1f: out <= 12'h222;
      20'h07f20: out <= 12'h000;
      20'h07f21: out <= 12'h660;
      20'h07f22: out <= 12'hbb0;
      20'h07f23: out <= 12'hee9;
      20'h07f24: out <= 12'hbb0;
      20'h07f25: out <= 12'hbb0;
      20'h07f26: out <= 12'h660;
      20'h07f27: out <= 12'h660;
      20'h07f28: out <= 12'h660;
      20'h07f29: out <= 12'h660;
      20'h07f2a: out <= 12'h660;
      20'h07f2b: out <= 12'h660;
      20'h07f2c: out <= 12'hee9;
      20'h07f2d: out <= 12'hbb0;
      20'h07f2e: out <= 12'h660;
      20'h07f2f: out <= 12'h000;
      20'h07f30: out <= 12'h222;
      20'h07f31: out <= 12'h660;
      20'h07f32: out <= 12'hbb0;
      20'h07f33: out <= 12'hee9;
      20'h07f34: out <= 12'hbb0;
      20'h07f35: out <= 12'h660;
      20'h07f36: out <= 12'h660;
      20'h07f37: out <= 12'h660;
      20'h07f38: out <= 12'h660;
      20'h07f39: out <= 12'h660;
      20'h07f3a: out <= 12'h660;
      20'h07f3b: out <= 12'h660;
      20'h07f3c: out <= 12'hee9;
      20'h07f3d: out <= 12'hbb0;
      20'h07f3e: out <= 12'h660;
      20'h07f3f: out <= 12'h222;
      20'h07f40: out <= 12'h000;
      20'h07f41: out <= 12'h000;
      20'h07f42: out <= 12'h660;
      20'h07f43: out <= 12'hee9;
      20'h07f44: out <= 12'hbb0;
      20'h07f45: out <= 12'h660;
      20'h07f46: out <= 12'h660;
      20'h07f47: out <= 12'h660;
      20'h07f48: out <= 12'h660;
      20'h07f49: out <= 12'h660;
      20'h07f4a: out <= 12'h660;
      20'h07f4b: out <= 12'h660;
      20'h07f4c: out <= 12'hbb0;
      20'h07f4d: out <= 12'hee9;
      20'h07f4e: out <= 12'h660;
      20'h07f4f: out <= 12'h000;
      20'h07f50: out <= 12'h222;
      20'h07f51: out <= 12'h222;
      20'h07f52: out <= 12'h660;
      20'h07f53: out <= 12'h660;
      20'h07f54: out <= 12'hbb0;
      20'h07f55: out <= 12'h660;
      20'h07f56: out <= 12'h660;
      20'h07f57: out <= 12'h660;
      20'h07f58: out <= 12'h660;
      20'h07f59: out <= 12'h660;
      20'h07f5a: out <= 12'h660;
      20'h07f5b: out <= 12'h660;
      20'h07f5c: out <= 12'hbb0;
      20'h07f5d: out <= 12'h660;
      20'h07f5e: out <= 12'h660;
      20'h07f5f: out <= 12'h222;
      20'h07f60: out <= 12'h603;
      20'h07f61: out <= 12'h603;
      20'h07f62: out <= 12'h603;
      20'h07f63: out <= 12'h603;
      20'h07f64: out <= 12'h603;
      20'h07f65: out <= 12'h603;
      20'h07f66: out <= 12'h603;
      20'h07f67: out <= 12'h603;
      20'h07f68: out <= 12'h603;
      20'h07f69: out <= 12'h603;
      20'h07f6a: out <= 12'h603;
      20'h07f6b: out <= 12'h603;
      20'h07f6c: out <= 12'hee9;
      20'h07f6d: out <= 12'hf87;
      20'h07f6e: out <= 12'hee9;
      20'h07f6f: out <= 12'hf87;
      20'h07f70: out <= 12'hf87;
      20'h07f71: out <= 12'hb27;
      20'h07f72: out <= 12'hf87;
      20'h07f73: out <= 12'hb27;
      20'h07f74: out <= 12'h603;
      20'h07f75: out <= 12'h603;
      20'h07f76: out <= 12'h603;
      20'h07f77: out <= 12'h603;
      20'h07f78: out <= 12'h603;
      20'h07f79: out <= 12'h603;
      20'h07f7a: out <= 12'h603;
      20'h07f7b: out <= 12'h603;
      20'h07f7c: out <= 12'h603;
      20'h07f7d: out <= 12'h603;
      20'h07f7e: out <= 12'h603;
      20'h07f7f: out <= 12'h603;
      20'h07f80: out <= 12'h603;
      20'h07f81: out <= 12'h603;
      20'h07f82: out <= 12'h603;
      20'h07f83: out <= 12'h603;
      20'h07f84: out <= 12'hee9;
      20'h07f85: out <= 12'hf87;
      20'h07f86: out <= 12'hee9;
      20'h07f87: out <= 12'hf87;
      20'h07f88: out <= 12'hf87;
      20'h07f89: out <= 12'hb27;
      20'h07f8a: out <= 12'hf87;
      20'h07f8b: out <= 12'hb27;
      20'h07f8c: out <= 12'h603;
      20'h07f8d: out <= 12'h603;
      20'h07f8e: out <= 12'h603;
      20'h07f8f: out <= 12'h603;
      20'h07f90: out <= 12'h603;
      20'h07f91: out <= 12'h603;
      20'h07f92: out <= 12'h603;
      20'h07f93: out <= 12'h603;
      20'h07f94: out <= 12'h603;
      20'h07f95: out <= 12'h603;
      20'h07f96: out <= 12'h603;
      20'h07f97: out <= 12'h603;
      20'h07f98: out <= 12'h603;
      20'h07f99: out <= 12'h603;
      20'h07f9a: out <= 12'h603;
      20'h07f9b: out <= 12'h603;
      20'h07f9c: out <= 12'h603;
      20'h07f9d: out <= 12'h603;
      20'h07f9e: out <= 12'h603;
      20'h07f9f: out <= 12'h603;
      20'h07fa0: out <= 12'h603;
      20'h07fa1: out <= 12'h603;
      20'h07fa2: out <= 12'h603;
      20'h07fa3: out <= 12'h603;
      20'h07fa4: out <= 12'h603;
      20'h07fa5: out <= 12'h603;
      20'h07fa6: out <= 12'h603;
      20'h07fa7: out <= 12'h603;
      20'h07fa8: out <= 12'h603;
      20'h07fa9: out <= 12'h603;
      20'h07faa: out <= 12'h603;
      20'h07fab: out <= 12'h603;
      20'h07fac: out <= 12'h603;
      20'h07fad: out <= 12'h603;
      20'h07fae: out <= 12'h603;
      20'h07faf: out <= 12'h603;
      20'h07fb0: out <= 12'h603;
      20'h07fb1: out <= 12'h603;
      20'h07fb2: out <= 12'h603;
      20'h07fb3: out <= 12'h603;
      20'h07fb4: out <= 12'h603;
      20'h07fb5: out <= 12'h603;
      20'h07fb6: out <= 12'h603;
      20'h07fb7: out <= 12'h603;
      20'h07fb8: out <= 12'hee9;
      20'h07fb9: out <= 12'hf87;
      20'h07fba: out <= 12'hee9;
      20'h07fbb: out <= 12'hf87;
      20'h07fbc: out <= 12'hf87;
      20'h07fbd: out <= 12'hb27;
      20'h07fbe: out <= 12'hf87;
      20'h07fbf: out <= 12'hb27;
      20'h07fc0: out <= 12'hee9;
      20'h07fc1: out <= 12'hf87;
      20'h07fc2: out <= 12'hee9;
      20'h07fc3: out <= 12'hf87;
      20'h07fc4: out <= 12'hf87;
      20'h07fc5: out <= 12'hb27;
      20'h07fc6: out <= 12'hf87;
      20'h07fc7: out <= 12'hb27;
      20'h07fc8: out <= 12'hee9;
      20'h07fc9: out <= 12'hf87;
      20'h07fca: out <= 12'hee9;
      20'h07fcb: out <= 12'hf87;
      20'h07fcc: out <= 12'hf87;
      20'h07fcd: out <= 12'hb27;
      20'h07fce: out <= 12'hf87;
      20'h07fcf: out <= 12'hb27;
      20'h07fd0: out <= 12'hee9;
      20'h07fd1: out <= 12'hf87;
      20'h07fd2: out <= 12'hee9;
      20'h07fd3: out <= 12'hf87;
      20'h07fd4: out <= 12'hf87;
      20'h07fd5: out <= 12'hb27;
      20'h07fd6: out <= 12'hf87;
      20'h07fd7: out <= 12'hb27;
      20'h07fd8: out <= 12'hee9;
      20'h07fd9: out <= 12'hf87;
      20'h07fda: out <= 12'hee9;
      20'h07fdb: out <= 12'hf87;
      20'h07fdc: out <= 12'hf87;
      20'h07fdd: out <= 12'hb27;
      20'h07fde: out <= 12'hf87;
      20'h07fdf: out <= 12'hb27;
      20'h07fe0: out <= 12'hee9;
      20'h07fe1: out <= 12'hf87;
      20'h07fe2: out <= 12'hee9;
      20'h07fe3: out <= 12'hf87;
      20'h07fe4: out <= 12'hf87;
      20'h07fe5: out <= 12'hb27;
      20'h07fe6: out <= 12'hf87;
      20'h07fe7: out <= 12'hb27;
      20'h07fe8: out <= 12'hee9;
      20'h07fe9: out <= 12'hf87;
      20'h07fea: out <= 12'hee9;
      20'h07feb: out <= 12'hf87;
      20'h07fec: out <= 12'hf87;
      20'h07fed: out <= 12'hb27;
      20'h07fee: out <= 12'hf87;
      20'h07fef: out <= 12'hb27;
      20'h07ff0: out <= 12'hee9;
      20'h07ff1: out <= 12'hf87;
      20'h07ff2: out <= 12'hee9;
      20'h07ff3: out <= 12'hf87;
      20'h07ff4: out <= 12'hf87;
      20'h07ff5: out <= 12'hb27;
      20'h07ff6: out <= 12'hf87;
      20'h07ff7: out <= 12'hb27;
      20'h07ff8: out <= 12'h000;
      20'h07ff9: out <= 12'hbb0;
      20'h07ffa: out <= 12'hee9;
      20'h07ffb: out <= 12'hbb0;
      20'h07ffc: out <= 12'h660;
      20'h07ffd: out <= 12'h660;
      20'h07ffe: out <= 12'hbb0;
      20'h07fff: out <= 12'hbb0;
      20'h08000: out <= 12'hee9;
      20'h08001: out <= 12'hee9;
      20'h08002: out <= 12'h660;
      20'h08003: out <= 12'h660;
      20'h08004: out <= 12'h660;
      20'h08005: out <= 12'hee9;
      20'h08006: out <= 12'hbb0;
      20'h08007: out <= 12'h000;
      20'h08008: out <= 12'h222;
      20'h08009: out <= 12'hbb0;
      20'h0800a: out <= 12'hee9;
      20'h0800b: out <= 12'hbb0;
      20'h0800c: out <= 12'h660;
      20'h0800d: out <= 12'h660;
      20'h0800e: out <= 12'hbb0;
      20'h0800f: out <= 12'hbb0;
      20'h08010: out <= 12'hee9;
      20'h08011: out <= 12'hee9;
      20'h08012: out <= 12'h660;
      20'h08013: out <= 12'h660;
      20'h08014: out <= 12'h660;
      20'h08015: out <= 12'hee9;
      20'h08016: out <= 12'hbb0;
      20'h08017: out <= 12'h222;
      20'h08018: out <= 12'h000;
      20'h08019: out <= 12'h000;
      20'h0801a: out <= 12'h660;
      20'h0801b: out <= 12'hee9;
      20'h0801c: out <= 12'hbb0;
      20'h0801d: out <= 12'hbb0;
      20'h0801e: out <= 12'h660;
      20'h0801f: out <= 12'h660;
      20'h08020: out <= 12'h660;
      20'h08021: out <= 12'h660;
      20'h08022: out <= 12'h660;
      20'h08023: out <= 12'hbb0;
      20'h08024: out <= 12'hbb0;
      20'h08025: out <= 12'hee9;
      20'h08026: out <= 12'h660;
      20'h08027: out <= 12'h000;
      20'h08028: out <= 12'h222;
      20'h08029: out <= 12'h222;
      20'h0802a: out <= 12'h660;
      20'h0802b: out <= 12'h660;
      20'h0802c: out <= 12'hbb0;
      20'h0802d: out <= 12'h660;
      20'h0802e: out <= 12'h660;
      20'h0802f: out <= 12'h660;
      20'h08030: out <= 12'h660;
      20'h08031: out <= 12'h660;
      20'h08032: out <= 12'h660;
      20'h08033: out <= 12'h660;
      20'h08034: out <= 12'hbb0;
      20'h08035: out <= 12'h660;
      20'h08036: out <= 12'h660;
      20'h08037: out <= 12'h222;
      20'h08038: out <= 12'h000;
      20'h08039: out <= 12'hbb0;
      20'h0803a: out <= 12'hee9;
      20'h0803b: out <= 12'h660;
      20'h0803c: out <= 12'h660;
      20'h0803d: out <= 12'h660;
      20'h0803e: out <= 12'hee9;
      20'h0803f: out <= 12'hee9;
      20'h08040: out <= 12'hbb0;
      20'h08041: out <= 12'hbb0;
      20'h08042: out <= 12'h660;
      20'h08043: out <= 12'h660;
      20'h08044: out <= 12'hbb0;
      20'h08045: out <= 12'hee9;
      20'h08046: out <= 12'hbb0;
      20'h08047: out <= 12'h000;
      20'h08048: out <= 12'h222;
      20'h08049: out <= 12'hbb0;
      20'h0804a: out <= 12'hee9;
      20'h0804b: out <= 12'h660;
      20'h0804c: out <= 12'h660;
      20'h0804d: out <= 12'h660;
      20'h0804e: out <= 12'hee9;
      20'h0804f: out <= 12'hee9;
      20'h08050: out <= 12'hbb0;
      20'h08051: out <= 12'hbb0;
      20'h08052: out <= 12'h660;
      20'h08053: out <= 12'h660;
      20'h08054: out <= 12'hbb0;
      20'h08055: out <= 12'hee9;
      20'h08056: out <= 12'hbb0;
      20'h08057: out <= 12'h222;
      20'h08058: out <= 12'h000;
      20'h08059: out <= 12'h000;
      20'h0805a: out <= 12'h660;
      20'h0805b: out <= 12'h660;
      20'h0805c: out <= 12'hbb0;
      20'h0805d: out <= 12'h660;
      20'h0805e: out <= 12'h660;
      20'h0805f: out <= 12'h660;
      20'h08060: out <= 12'h660;
      20'h08061: out <= 12'h660;
      20'h08062: out <= 12'h660;
      20'h08063: out <= 12'h660;
      20'h08064: out <= 12'hbb0;
      20'h08065: out <= 12'h660;
      20'h08066: out <= 12'h660;
      20'h08067: out <= 12'h000;
      20'h08068: out <= 12'h222;
      20'h08069: out <= 12'h222;
      20'h0806a: out <= 12'h660;
      20'h0806b: out <= 12'hee9;
      20'h0806c: out <= 12'hbb0;
      20'h0806d: out <= 12'h660;
      20'h0806e: out <= 12'h660;
      20'h0806f: out <= 12'h660;
      20'h08070: out <= 12'h660;
      20'h08071: out <= 12'h660;
      20'h08072: out <= 12'h660;
      20'h08073: out <= 12'h660;
      20'h08074: out <= 12'hbb0;
      20'h08075: out <= 12'hee9;
      20'h08076: out <= 12'h660;
      20'h08077: out <= 12'h222;
      20'h08078: out <= 12'h603;
      20'h08079: out <= 12'h603;
      20'h0807a: out <= 12'h603;
      20'h0807b: out <= 12'h603;
      20'h0807c: out <= 12'h603;
      20'h0807d: out <= 12'h603;
      20'h0807e: out <= 12'h603;
      20'h0807f: out <= 12'h603;
      20'h08080: out <= 12'h603;
      20'h08081: out <= 12'h603;
      20'h08082: out <= 12'h603;
      20'h08083: out <= 12'h603;
      20'h08084: out <= 12'hee9;
      20'h08085: out <= 12'hf87;
      20'h08086: out <= 12'hee9;
      20'h08087: out <= 12'hb27;
      20'h08088: out <= 12'hb27;
      20'h08089: out <= 12'hb27;
      20'h0808a: out <= 12'hf87;
      20'h0808b: out <= 12'hb27;
      20'h0808c: out <= 12'h603;
      20'h0808d: out <= 12'h603;
      20'h0808e: out <= 12'h603;
      20'h0808f: out <= 12'h603;
      20'h08090: out <= 12'h603;
      20'h08091: out <= 12'h603;
      20'h08092: out <= 12'h603;
      20'h08093: out <= 12'h603;
      20'h08094: out <= 12'h603;
      20'h08095: out <= 12'h603;
      20'h08096: out <= 12'h603;
      20'h08097: out <= 12'h603;
      20'h08098: out <= 12'h603;
      20'h08099: out <= 12'h603;
      20'h0809a: out <= 12'h603;
      20'h0809b: out <= 12'h603;
      20'h0809c: out <= 12'hee9;
      20'h0809d: out <= 12'hf87;
      20'h0809e: out <= 12'hee9;
      20'h0809f: out <= 12'hb27;
      20'h080a0: out <= 12'hb27;
      20'h080a1: out <= 12'hb27;
      20'h080a2: out <= 12'hf87;
      20'h080a3: out <= 12'hb27;
      20'h080a4: out <= 12'h603;
      20'h080a5: out <= 12'h603;
      20'h080a6: out <= 12'h603;
      20'h080a7: out <= 12'h603;
      20'h080a8: out <= 12'h603;
      20'h080a9: out <= 12'h603;
      20'h080aa: out <= 12'h603;
      20'h080ab: out <= 12'h603;
      20'h080ac: out <= 12'h603;
      20'h080ad: out <= 12'h603;
      20'h080ae: out <= 12'h603;
      20'h080af: out <= 12'h603;
      20'h080b0: out <= 12'h603;
      20'h080b1: out <= 12'h603;
      20'h080b2: out <= 12'h603;
      20'h080b3: out <= 12'h603;
      20'h080b4: out <= 12'h603;
      20'h080b5: out <= 12'h603;
      20'h080b6: out <= 12'h603;
      20'h080b7: out <= 12'h603;
      20'h080b8: out <= 12'h603;
      20'h080b9: out <= 12'h603;
      20'h080ba: out <= 12'h603;
      20'h080bb: out <= 12'h603;
      20'h080bc: out <= 12'h603;
      20'h080bd: out <= 12'h603;
      20'h080be: out <= 12'h603;
      20'h080bf: out <= 12'h603;
      20'h080c0: out <= 12'h603;
      20'h080c1: out <= 12'h603;
      20'h080c2: out <= 12'h603;
      20'h080c3: out <= 12'h603;
      20'h080c4: out <= 12'h603;
      20'h080c5: out <= 12'h603;
      20'h080c6: out <= 12'h603;
      20'h080c7: out <= 12'h603;
      20'h080c8: out <= 12'h603;
      20'h080c9: out <= 12'h603;
      20'h080ca: out <= 12'h603;
      20'h080cb: out <= 12'h603;
      20'h080cc: out <= 12'h603;
      20'h080cd: out <= 12'h603;
      20'h080ce: out <= 12'h603;
      20'h080cf: out <= 12'h603;
      20'h080d0: out <= 12'hee9;
      20'h080d1: out <= 12'hf87;
      20'h080d2: out <= 12'hee9;
      20'h080d3: out <= 12'hb27;
      20'h080d4: out <= 12'hb27;
      20'h080d5: out <= 12'hb27;
      20'h080d6: out <= 12'hf87;
      20'h080d7: out <= 12'hb27;
      20'h080d8: out <= 12'hee9;
      20'h080d9: out <= 12'hf87;
      20'h080da: out <= 12'hee9;
      20'h080db: out <= 12'hb27;
      20'h080dc: out <= 12'hb27;
      20'h080dd: out <= 12'hb27;
      20'h080de: out <= 12'hf87;
      20'h080df: out <= 12'hb27;
      20'h080e0: out <= 12'hee9;
      20'h080e1: out <= 12'hf87;
      20'h080e2: out <= 12'hee9;
      20'h080e3: out <= 12'hb27;
      20'h080e4: out <= 12'hb27;
      20'h080e5: out <= 12'hb27;
      20'h080e6: out <= 12'hf87;
      20'h080e7: out <= 12'hb27;
      20'h080e8: out <= 12'hee9;
      20'h080e9: out <= 12'hf87;
      20'h080ea: out <= 12'hee9;
      20'h080eb: out <= 12'hb27;
      20'h080ec: out <= 12'hb27;
      20'h080ed: out <= 12'hb27;
      20'h080ee: out <= 12'hf87;
      20'h080ef: out <= 12'hb27;
      20'h080f0: out <= 12'hee9;
      20'h080f1: out <= 12'hf87;
      20'h080f2: out <= 12'hee9;
      20'h080f3: out <= 12'hb27;
      20'h080f4: out <= 12'hb27;
      20'h080f5: out <= 12'hb27;
      20'h080f6: out <= 12'hf87;
      20'h080f7: out <= 12'hb27;
      20'h080f8: out <= 12'hee9;
      20'h080f9: out <= 12'hf87;
      20'h080fa: out <= 12'hee9;
      20'h080fb: out <= 12'hb27;
      20'h080fc: out <= 12'hb27;
      20'h080fd: out <= 12'hb27;
      20'h080fe: out <= 12'hf87;
      20'h080ff: out <= 12'hb27;
      20'h08100: out <= 12'hee9;
      20'h08101: out <= 12'hf87;
      20'h08102: out <= 12'hee9;
      20'h08103: out <= 12'hb27;
      20'h08104: out <= 12'hb27;
      20'h08105: out <= 12'hb27;
      20'h08106: out <= 12'hf87;
      20'h08107: out <= 12'hb27;
      20'h08108: out <= 12'hee9;
      20'h08109: out <= 12'hf87;
      20'h0810a: out <= 12'hee9;
      20'h0810b: out <= 12'hb27;
      20'h0810c: out <= 12'hb27;
      20'h0810d: out <= 12'hb27;
      20'h0810e: out <= 12'hf87;
      20'h0810f: out <= 12'hb27;
      20'h08110: out <= 12'h000;
      20'h08111: out <= 12'hbb0;
      20'h08112: out <= 12'hee9;
      20'h08113: out <= 12'hbb0;
      20'h08114: out <= 12'h660;
      20'h08115: out <= 12'h660;
      20'h08116: out <= 12'hbb0;
      20'h08117: out <= 12'hbb0;
      20'h08118: out <= 12'hee9;
      20'h08119: out <= 12'hee9;
      20'h0811a: out <= 12'h660;
      20'h0811b: out <= 12'hbb0;
      20'h0811c: out <= 12'h660;
      20'h0811d: out <= 12'h660;
      20'h0811e: out <= 12'h660;
      20'h0811f: out <= 12'h660;
      20'h08120: out <= 12'h222;
      20'h08121: out <= 12'hbb0;
      20'h08122: out <= 12'hee9;
      20'h08123: out <= 12'hbb0;
      20'h08124: out <= 12'h660;
      20'h08125: out <= 12'h660;
      20'h08126: out <= 12'hbb0;
      20'h08127: out <= 12'hbb0;
      20'h08128: out <= 12'hee9;
      20'h08129: out <= 12'hee9;
      20'h0812a: out <= 12'h660;
      20'h0812b: out <= 12'hbb0;
      20'h0812c: out <= 12'h660;
      20'h0812d: out <= 12'h660;
      20'h0812e: out <= 12'h660;
      20'h0812f: out <= 12'h660;
      20'h08130: out <= 12'h000;
      20'h08131: out <= 12'h000;
      20'h08132: out <= 12'h660;
      20'h08133: out <= 12'h660;
      20'h08134: out <= 12'hbb0;
      20'h08135: out <= 12'h660;
      20'h08136: out <= 12'hee9;
      20'h08137: out <= 12'hee9;
      20'h08138: out <= 12'hee9;
      20'h08139: out <= 12'hee9;
      20'h0813a: out <= 12'hee9;
      20'h0813b: out <= 12'h660;
      20'h0813c: out <= 12'hbb0;
      20'h0813d: out <= 12'h660;
      20'h0813e: out <= 12'h660;
      20'h0813f: out <= 12'h000;
      20'h08140: out <= 12'h222;
      20'h08141: out <= 12'h222;
      20'h08142: out <= 12'h660;
      20'h08143: out <= 12'hee9;
      20'h08144: out <= 12'hbb0;
      20'h08145: out <= 12'h660;
      20'h08146: out <= 12'hee9;
      20'h08147: out <= 12'hee9;
      20'h08148: out <= 12'hee9;
      20'h08149: out <= 12'hee9;
      20'h0814a: out <= 12'hee9;
      20'h0814b: out <= 12'h660;
      20'h0814c: out <= 12'hbb0;
      20'h0814d: out <= 12'hee9;
      20'h0814e: out <= 12'h660;
      20'h0814f: out <= 12'h222;
      20'h08150: out <= 12'h660;
      20'h08151: out <= 12'h660;
      20'h08152: out <= 12'h660;
      20'h08153: out <= 12'h660;
      20'h08154: out <= 12'hbb0;
      20'h08155: out <= 12'h660;
      20'h08156: out <= 12'hee9;
      20'h08157: out <= 12'hee9;
      20'h08158: out <= 12'hbb0;
      20'h08159: out <= 12'hbb0;
      20'h0815a: out <= 12'h660;
      20'h0815b: out <= 12'h660;
      20'h0815c: out <= 12'hbb0;
      20'h0815d: out <= 12'hee9;
      20'h0815e: out <= 12'hbb0;
      20'h0815f: out <= 12'h000;
      20'h08160: out <= 12'h660;
      20'h08161: out <= 12'h660;
      20'h08162: out <= 12'h660;
      20'h08163: out <= 12'h660;
      20'h08164: out <= 12'hbb0;
      20'h08165: out <= 12'h660;
      20'h08166: out <= 12'hee9;
      20'h08167: out <= 12'hee9;
      20'h08168: out <= 12'hbb0;
      20'h08169: out <= 12'hbb0;
      20'h0816a: out <= 12'h660;
      20'h0816b: out <= 12'h660;
      20'h0816c: out <= 12'hbb0;
      20'h0816d: out <= 12'hee9;
      20'h0816e: out <= 12'hbb0;
      20'h0816f: out <= 12'h222;
      20'h08170: out <= 12'h000;
      20'h08171: out <= 12'h000;
      20'h08172: out <= 12'h660;
      20'h08173: out <= 12'hee9;
      20'h08174: out <= 12'hbb0;
      20'h08175: out <= 12'h660;
      20'h08176: out <= 12'hbb0;
      20'h08177: out <= 12'hbb0;
      20'h08178: out <= 12'hbb0;
      20'h08179: out <= 12'hbb0;
      20'h0817a: out <= 12'hbb0;
      20'h0817b: out <= 12'h660;
      20'h0817c: out <= 12'hbb0;
      20'h0817d: out <= 12'hee9;
      20'h0817e: out <= 12'h660;
      20'h0817f: out <= 12'h000;
      20'h08180: out <= 12'h222;
      20'h08181: out <= 12'h222;
      20'h08182: out <= 12'h660;
      20'h08183: out <= 12'h660;
      20'h08184: out <= 12'hbb0;
      20'h08185: out <= 12'h660;
      20'h08186: out <= 12'hbb0;
      20'h08187: out <= 12'hbb0;
      20'h08188: out <= 12'hbb0;
      20'h08189: out <= 12'hbb0;
      20'h0818a: out <= 12'hbb0;
      20'h0818b: out <= 12'h660;
      20'h0818c: out <= 12'hbb0;
      20'h0818d: out <= 12'h660;
      20'h0818e: out <= 12'h660;
      20'h0818f: out <= 12'h222;
      20'h08190: out <= 12'h603;
      20'h08191: out <= 12'h603;
      20'h08192: out <= 12'h603;
      20'h08193: out <= 12'h603;
      20'h08194: out <= 12'h603;
      20'h08195: out <= 12'h603;
      20'h08196: out <= 12'h603;
      20'h08197: out <= 12'h603;
      20'h08198: out <= 12'h603;
      20'h08199: out <= 12'h603;
      20'h0819a: out <= 12'h603;
      20'h0819b: out <= 12'h603;
      20'h0819c: out <= 12'hee9;
      20'h0819d: out <= 12'hf87;
      20'h0819e: out <= 12'hf87;
      20'h0819f: out <= 12'hf87;
      20'h081a0: out <= 12'hf87;
      20'h081a1: out <= 12'hf87;
      20'h081a2: out <= 12'hf87;
      20'h081a3: out <= 12'hb27;
      20'h081a4: out <= 12'h603;
      20'h081a5: out <= 12'h603;
      20'h081a6: out <= 12'h603;
      20'h081a7: out <= 12'h603;
      20'h081a8: out <= 12'h603;
      20'h081a9: out <= 12'h603;
      20'h081aa: out <= 12'h603;
      20'h081ab: out <= 12'h603;
      20'h081ac: out <= 12'h603;
      20'h081ad: out <= 12'h603;
      20'h081ae: out <= 12'h603;
      20'h081af: out <= 12'h603;
      20'h081b0: out <= 12'h603;
      20'h081b1: out <= 12'h603;
      20'h081b2: out <= 12'h603;
      20'h081b3: out <= 12'h603;
      20'h081b4: out <= 12'hee9;
      20'h081b5: out <= 12'hf87;
      20'h081b6: out <= 12'hf87;
      20'h081b7: out <= 12'hf87;
      20'h081b8: out <= 12'hf87;
      20'h081b9: out <= 12'hf87;
      20'h081ba: out <= 12'hf87;
      20'h081bb: out <= 12'hb27;
      20'h081bc: out <= 12'h603;
      20'h081bd: out <= 12'h603;
      20'h081be: out <= 12'h603;
      20'h081bf: out <= 12'h603;
      20'h081c0: out <= 12'h603;
      20'h081c1: out <= 12'h603;
      20'h081c2: out <= 12'h603;
      20'h081c3: out <= 12'h603;
      20'h081c4: out <= 12'h603;
      20'h081c5: out <= 12'h603;
      20'h081c6: out <= 12'h603;
      20'h081c7: out <= 12'h603;
      20'h081c8: out <= 12'h603;
      20'h081c9: out <= 12'h603;
      20'h081ca: out <= 12'h603;
      20'h081cb: out <= 12'h603;
      20'h081cc: out <= 12'h603;
      20'h081cd: out <= 12'h603;
      20'h081ce: out <= 12'h603;
      20'h081cf: out <= 12'h603;
      20'h081d0: out <= 12'h603;
      20'h081d1: out <= 12'h603;
      20'h081d2: out <= 12'h603;
      20'h081d3: out <= 12'h603;
      20'h081d4: out <= 12'h603;
      20'h081d5: out <= 12'h603;
      20'h081d6: out <= 12'h603;
      20'h081d7: out <= 12'h603;
      20'h081d8: out <= 12'h603;
      20'h081d9: out <= 12'h603;
      20'h081da: out <= 12'h603;
      20'h081db: out <= 12'h603;
      20'h081dc: out <= 12'h603;
      20'h081dd: out <= 12'h603;
      20'h081de: out <= 12'h603;
      20'h081df: out <= 12'h603;
      20'h081e0: out <= 12'h603;
      20'h081e1: out <= 12'h603;
      20'h081e2: out <= 12'h603;
      20'h081e3: out <= 12'h603;
      20'h081e4: out <= 12'h603;
      20'h081e5: out <= 12'h603;
      20'h081e6: out <= 12'h603;
      20'h081e7: out <= 12'h603;
      20'h081e8: out <= 12'hee9;
      20'h081e9: out <= 12'hf87;
      20'h081ea: out <= 12'hf87;
      20'h081eb: out <= 12'hf87;
      20'h081ec: out <= 12'hf87;
      20'h081ed: out <= 12'hf87;
      20'h081ee: out <= 12'hf87;
      20'h081ef: out <= 12'hb27;
      20'h081f0: out <= 12'hee9;
      20'h081f1: out <= 12'hf87;
      20'h081f2: out <= 12'hf87;
      20'h081f3: out <= 12'hf87;
      20'h081f4: out <= 12'hf87;
      20'h081f5: out <= 12'hf87;
      20'h081f6: out <= 12'hf87;
      20'h081f7: out <= 12'hb27;
      20'h081f8: out <= 12'hee9;
      20'h081f9: out <= 12'hf87;
      20'h081fa: out <= 12'hf87;
      20'h081fb: out <= 12'hf87;
      20'h081fc: out <= 12'hf87;
      20'h081fd: out <= 12'hf87;
      20'h081fe: out <= 12'hf87;
      20'h081ff: out <= 12'hb27;
      20'h08200: out <= 12'hee9;
      20'h08201: out <= 12'hf87;
      20'h08202: out <= 12'hf87;
      20'h08203: out <= 12'hf87;
      20'h08204: out <= 12'hf87;
      20'h08205: out <= 12'hf87;
      20'h08206: out <= 12'hf87;
      20'h08207: out <= 12'hb27;
      20'h08208: out <= 12'hee9;
      20'h08209: out <= 12'hf87;
      20'h0820a: out <= 12'hf87;
      20'h0820b: out <= 12'hf87;
      20'h0820c: out <= 12'hf87;
      20'h0820d: out <= 12'hf87;
      20'h0820e: out <= 12'hf87;
      20'h0820f: out <= 12'hb27;
      20'h08210: out <= 12'hee9;
      20'h08211: out <= 12'hf87;
      20'h08212: out <= 12'hf87;
      20'h08213: out <= 12'hf87;
      20'h08214: out <= 12'hf87;
      20'h08215: out <= 12'hf87;
      20'h08216: out <= 12'hf87;
      20'h08217: out <= 12'hb27;
      20'h08218: out <= 12'hee9;
      20'h08219: out <= 12'hf87;
      20'h0821a: out <= 12'hf87;
      20'h0821b: out <= 12'hf87;
      20'h0821c: out <= 12'hf87;
      20'h0821d: out <= 12'hf87;
      20'h0821e: out <= 12'hf87;
      20'h0821f: out <= 12'hb27;
      20'h08220: out <= 12'hee9;
      20'h08221: out <= 12'hf87;
      20'h08222: out <= 12'hf87;
      20'h08223: out <= 12'hf87;
      20'h08224: out <= 12'hf87;
      20'h08225: out <= 12'hf87;
      20'h08226: out <= 12'hf87;
      20'h08227: out <= 12'hb27;
      20'h08228: out <= 12'h000;
      20'h08229: out <= 12'hbb0;
      20'h0822a: out <= 12'hee9;
      20'h0822b: out <= 12'hbb0;
      20'h0822c: out <= 12'h660;
      20'h0822d: out <= 12'h660;
      20'h0822e: out <= 12'hbb0;
      20'h0822f: out <= 12'hbb0;
      20'h08230: out <= 12'hee9;
      20'h08231: out <= 12'hee9;
      20'h08232: out <= 12'h660;
      20'h08233: out <= 12'hee9;
      20'h08234: out <= 12'hee9;
      20'h08235: out <= 12'hee9;
      20'h08236: out <= 12'hee9;
      20'h08237: out <= 12'hee9;
      20'h08238: out <= 12'h222;
      20'h08239: out <= 12'hbb0;
      20'h0823a: out <= 12'hee9;
      20'h0823b: out <= 12'hbb0;
      20'h0823c: out <= 12'h660;
      20'h0823d: out <= 12'h660;
      20'h0823e: out <= 12'hbb0;
      20'h0823f: out <= 12'hbb0;
      20'h08240: out <= 12'hee9;
      20'h08241: out <= 12'hee9;
      20'h08242: out <= 12'h660;
      20'h08243: out <= 12'hee9;
      20'h08244: out <= 12'hee9;
      20'h08245: out <= 12'hee9;
      20'h08246: out <= 12'hee9;
      20'h08247: out <= 12'hee9;
      20'h08248: out <= 12'h000;
      20'h08249: out <= 12'h000;
      20'h0824a: out <= 12'h660;
      20'h0824b: out <= 12'hee9;
      20'h0824c: out <= 12'hbb0;
      20'h0824d: out <= 12'h660;
      20'h0824e: out <= 12'hee9;
      20'h0824f: out <= 12'hee9;
      20'h08250: out <= 12'hee9;
      20'h08251: out <= 12'hee9;
      20'h08252: out <= 12'hee9;
      20'h08253: out <= 12'h660;
      20'h08254: out <= 12'hbb0;
      20'h08255: out <= 12'hee9;
      20'h08256: out <= 12'h660;
      20'h08257: out <= 12'h000;
      20'h08258: out <= 12'h222;
      20'h08259: out <= 12'h222;
      20'h0825a: out <= 12'h660;
      20'h0825b: out <= 12'h660;
      20'h0825c: out <= 12'hbb0;
      20'h0825d: out <= 12'h660;
      20'h0825e: out <= 12'hee9;
      20'h0825f: out <= 12'hee9;
      20'h08260: out <= 12'hee9;
      20'h08261: out <= 12'hee9;
      20'h08262: out <= 12'hee9;
      20'h08263: out <= 12'h660;
      20'h08264: out <= 12'hbb0;
      20'h08265: out <= 12'h660;
      20'h08266: out <= 12'h660;
      20'h08267: out <= 12'h222;
      20'h08268: out <= 12'hee9;
      20'h08269: out <= 12'hee9;
      20'h0826a: out <= 12'hee9;
      20'h0826b: out <= 12'hee9;
      20'h0826c: out <= 12'hee9;
      20'h0826d: out <= 12'h660;
      20'h0826e: out <= 12'hee9;
      20'h0826f: out <= 12'hee9;
      20'h08270: out <= 12'hbb0;
      20'h08271: out <= 12'hbb0;
      20'h08272: out <= 12'h660;
      20'h08273: out <= 12'h660;
      20'h08274: out <= 12'hbb0;
      20'h08275: out <= 12'hee9;
      20'h08276: out <= 12'hbb0;
      20'h08277: out <= 12'h000;
      20'h08278: out <= 12'hee9;
      20'h08279: out <= 12'hee9;
      20'h0827a: out <= 12'hee9;
      20'h0827b: out <= 12'hee9;
      20'h0827c: out <= 12'hee9;
      20'h0827d: out <= 12'h660;
      20'h0827e: out <= 12'hee9;
      20'h0827f: out <= 12'hee9;
      20'h08280: out <= 12'hbb0;
      20'h08281: out <= 12'hbb0;
      20'h08282: out <= 12'h660;
      20'h08283: out <= 12'h660;
      20'h08284: out <= 12'hbb0;
      20'h08285: out <= 12'hee9;
      20'h08286: out <= 12'hbb0;
      20'h08287: out <= 12'h222;
      20'h08288: out <= 12'h000;
      20'h08289: out <= 12'h000;
      20'h0828a: out <= 12'h660;
      20'h0828b: out <= 12'h660;
      20'h0828c: out <= 12'hbb0;
      20'h0828d: out <= 12'h660;
      20'h0828e: out <= 12'hbb0;
      20'h0828f: out <= 12'hbb0;
      20'h08290: out <= 12'hbb0;
      20'h08291: out <= 12'hbb0;
      20'h08292: out <= 12'hbb0;
      20'h08293: out <= 12'h660;
      20'h08294: out <= 12'hbb0;
      20'h08295: out <= 12'h660;
      20'h08296: out <= 12'h660;
      20'h08297: out <= 12'h000;
      20'h08298: out <= 12'h222;
      20'h08299: out <= 12'h222;
      20'h0829a: out <= 12'h660;
      20'h0829b: out <= 12'hee9;
      20'h0829c: out <= 12'hbb0;
      20'h0829d: out <= 12'h660;
      20'h0829e: out <= 12'hbb0;
      20'h0829f: out <= 12'hbb0;
      20'h082a0: out <= 12'hbb0;
      20'h082a1: out <= 12'hbb0;
      20'h082a2: out <= 12'hbb0;
      20'h082a3: out <= 12'h660;
      20'h082a4: out <= 12'hbb0;
      20'h082a5: out <= 12'hee9;
      20'h082a6: out <= 12'h660;
      20'h082a7: out <= 12'h222;
      20'h082a8: out <= 12'h603;
      20'h082a9: out <= 12'h603;
      20'h082aa: out <= 12'h603;
      20'h082ab: out <= 12'h603;
      20'h082ac: out <= 12'h603;
      20'h082ad: out <= 12'h603;
      20'h082ae: out <= 12'h603;
      20'h082af: out <= 12'h603;
      20'h082b0: out <= 12'h603;
      20'h082b1: out <= 12'h603;
      20'h082b2: out <= 12'h603;
      20'h082b3: out <= 12'h603;
      20'h082b4: out <= 12'hb27;
      20'h082b5: out <= 12'hb27;
      20'h082b6: out <= 12'hb27;
      20'h082b7: out <= 12'hb27;
      20'h082b8: out <= 12'hb27;
      20'h082b9: out <= 12'hb27;
      20'h082ba: out <= 12'hb27;
      20'h082bb: out <= 12'hb27;
      20'h082bc: out <= 12'h603;
      20'h082bd: out <= 12'h603;
      20'h082be: out <= 12'h603;
      20'h082bf: out <= 12'h603;
      20'h082c0: out <= 12'h603;
      20'h082c1: out <= 12'h603;
      20'h082c2: out <= 12'h603;
      20'h082c3: out <= 12'h603;
      20'h082c4: out <= 12'h603;
      20'h082c5: out <= 12'h603;
      20'h082c6: out <= 12'h603;
      20'h082c7: out <= 12'h603;
      20'h082c8: out <= 12'h603;
      20'h082c9: out <= 12'h603;
      20'h082ca: out <= 12'h603;
      20'h082cb: out <= 12'h603;
      20'h082cc: out <= 12'hb27;
      20'h082cd: out <= 12'hb27;
      20'h082ce: out <= 12'hb27;
      20'h082cf: out <= 12'hb27;
      20'h082d0: out <= 12'hb27;
      20'h082d1: out <= 12'hb27;
      20'h082d2: out <= 12'hb27;
      20'h082d3: out <= 12'hb27;
      20'h082d4: out <= 12'h603;
      20'h082d5: out <= 12'h603;
      20'h082d6: out <= 12'h603;
      20'h082d7: out <= 12'h603;
      20'h082d8: out <= 12'h603;
      20'h082d9: out <= 12'h603;
      20'h082da: out <= 12'h603;
      20'h082db: out <= 12'h603;
      20'h082dc: out <= 12'h603;
      20'h082dd: out <= 12'h603;
      20'h082de: out <= 12'h603;
      20'h082df: out <= 12'h603;
      20'h082e0: out <= 12'h603;
      20'h082e1: out <= 12'h603;
      20'h082e2: out <= 12'h603;
      20'h082e3: out <= 12'h603;
      20'h082e4: out <= 12'h603;
      20'h082e5: out <= 12'h603;
      20'h082e6: out <= 12'h603;
      20'h082e7: out <= 12'h603;
      20'h082e8: out <= 12'h603;
      20'h082e9: out <= 12'h603;
      20'h082ea: out <= 12'h603;
      20'h082eb: out <= 12'h603;
      20'h082ec: out <= 12'h603;
      20'h082ed: out <= 12'h603;
      20'h082ee: out <= 12'h603;
      20'h082ef: out <= 12'h603;
      20'h082f0: out <= 12'h603;
      20'h082f1: out <= 12'h603;
      20'h082f2: out <= 12'h603;
      20'h082f3: out <= 12'h603;
      20'h082f4: out <= 12'h603;
      20'h082f5: out <= 12'h603;
      20'h082f6: out <= 12'h603;
      20'h082f7: out <= 12'h603;
      20'h082f8: out <= 12'h603;
      20'h082f9: out <= 12'h603;
      20'h082fa: out <= 12'h603;
      20'h082fb: out <= 12'h603;
      20'h082fc: out <= 12'h603;
      20'h082fd: out <= 12'h603;
      20'h082fe: out <= 12'h603;
      20'h082ff: out <= 12'h603;
      20'h08300: out <= 12'hb27;
      20'h08301: out <= 12'hb27;
      20'h08302: out <= 12'hb27;
      20'h08303: out <= 12'hb27;
      20'h08304: out <= 12'hb27;
      20'h08305: out <= 12'hb27;
      20'h08306: out <= 12'hb27;
      20'h08307: out <= 12'hb27;
      20'h08308: out <= 12'hb27;
      20'h08309: out <= 12'hb27;
      20'h0830a: out <= 12'hb27;
      20'h0830b: out <= 12'hb27;
      20'h0830c: out <= 12'hb27;
      20'h0830d: out <= 12'hb27;
      20'h0830e: out <= 12'hb27;
      20'h0830f: out <= 12'hb27;
      20'h08310: out <= 12'hb27;
      20'h08311: out <= 12'hb27;
      20'h08312: out <= 12'hb27;
      20'h08313: out <= 12'hb27;
      20'h08314: out <= 12'hb27;
      20'h08315: out <= 12'hb27;
      20'h08316: out <= 12'hb27;
      20'h08317: out <= 12'hb27;
      20'h08318: out <= 12'hb27;
      20'h08319: out <= 12'hb27;
      20'h0831a: out <= 12'hb27;
      20'h0831b: out <= 12'hb27;
      20'h0831c: out <= 12'hb27;
      20'h0831d: out <= 12'hb27;
      20'h0831e: out <= 12'hb27;
      20'h0831f: out <= 12'hb27;
      20'h08320: out <= 12'hb27;
      20'h08321: out <= 12'hb27;
      20'h08322: out <= 12'hb27;
      20'h08323: out <= 12'hb27;
      20'h08324: out <= 12'hb27;
      20'h08325: out <= 12'hb27;
      20'h08326: out <= 12'hb27;
      20'h08327: out <= 12'hb27;
      20'h08328: out <= 12'hb27;
      20'h08329: out <= 12'hb27;
      20'h0832a: out <= 12'hb27;
      20'h0832b: out <= 12'hb27;
      20'h0832c: out <= 12'hb27;
      20'h0832d: out <= 12'hb27;
      20'h0832e: out <= 12'hb27;
      20'h0832f: out <= 12'hb27;
      20'h08330: out <= 12'hb27;
      20'h08331: out <= 12'hb27;
      20'h08332: out <= 12'hb27;
      20'h08333: out <= 12'hb27;
      20'h08334: out <= 12'hb27;
      20'h08335: out <= 12'hb27;
      20'h08336: out <= 12'hb27;
      20'h08337: out <= 12'hb27;
      20'h08338: out <= 12'hb27;
      20'h08339: out <= 12'hb27;
      20'h0833a: out <= 12'hb27;
      20'h0833b: out <= 12'hb27;
      20'h0833c: out <= 12'hb27;
      20'h0833d: out <= 12'hb27;
      20'h0833e: out <= 12'hb27;
      20'h0833f: out <= 12'hb27;
      20'h08340: out <= 12'h000;
      20'h08341: out <= 12'hbb0;
      20'h08342: out <= 12'hee9;
      20'h08343: out <= 12'hbb0;
      20'h08344: out <= 12'h660;
      20'h08345: out <= 12'h660;
      20'h08346: out <= 12'hbb0;
      20'h08347: out <= 12'hbb0;
      20'h08348: out <= 12'hee9;
      20'h08349: out <= 12'hee9;
      20'h0834a: out <= 12'h660;
      20'h0834b: out <= 12'hbb0;
      20'h0834c: out <= 12'h660;
      20'h0834d: out <= 12'h660;
      20'h0834e: out <= 12'h660;
      20'h0834f: out <= 12'h660;
      20'h08350: out <= 12'h222;
      20'h08351: out <= 12'hbb0;
      20'h08352: out <= 12'hee9;
      20'h08353: out <= 12'hbb0;
      20'h08354: out <= 12'h660;
      20'h08355: out <= 12'h660;
      20'h08356: out <= 12'hbb0;
      20'h08357: out <= 12'hbb0;
      20'h08358: out <= 12'hee9;
      20'h08359: out <= 12'hee9;
      20'h0835a: out <= 12'h660;
      20'h0835b: out <= 12'hbb0;
      20'h0835c: out <= 12'h660;
      20'h0835d: out <= 12'h660;
      20'h0835e: out <= 12'h660;
      20'h0835f: out <= 12'h660;
      20'h08360: out <= 12'h000;
      20'h08361: out <= 12'h000;
      20'h08362: out <= 12'h660;
      20'h08363: out <= 12'h660;
      20'h08364: out <= 12'hbb0;
      20'h08365: out <= 12'h660;
      20'h08366: out <= 12'hbb0;
      20'h08367: out <= 12'hbb0;
      20'h08368: out <= 12'hbb0;
      20'h08369: out <= 12'hbb0;
      20'h0836a: out <= 12'hbb0;
      20'h0836b: out <= 12'h660;
      20'h0836c: out <= 12'hbb0;
      20'h0836d: out <= 12'h660;
      20'h0836e: out <= 12'h660;
      20'h0836f: out <= 12'h000;
      20'h08370: out <= 12'h222;
      20'h08371: out <= 12'h222;
      20'h08372: out <= 12'h660;
      20'h08373: out <= 12'hee9;
      20'h08374: out <= 12'hbb0;
      20'h08375: out <= 12'h660;
      20'h08376: out <= 12'hbb0;
      20'h08377: out <= 12'hbb0;
      20'h08378: out <= 12'hbb0;
      20'h08379: out <= 12'hbb0;
      20'h0837a: out <= 12'hbb0;
      20'h0837b: out <= 12'h660;
      20'h0837c: out <= 12'hbb0;
      20'h0837d: out <= 12'hee9;
      20'h0837e: out <= 12'h660;
      20'h0837f: out <= 12'h222;
      20'h08380: out <= 12'h660;
      20'h08381: out <= 12'h660;
      20'h08382: out <= 12'h660;
      20'h08383: out <= 12'h660;
      20'h08384: out <= 12'hbb0;
      20'h08385: out <= 12'h660;
      20'h08386: out <= 12'hee9;
      20'h08387: out <= 12'hee9;
      20'h08388: out <= 12'hbb0;
      20'h08389: out <= 12'hbb0;
      20'h0838a: out <= 12'h660;
      20'h0838b: out <= 12'h660;
      20'h0838c: out <= 12'hbb0;
      20'h0838d: out <= 12'hee9;
      20'h0838e: out <= 12'hbb0;
      20'h0838f: out <= 12'h000;
      20'h08390: out <= 12'h660;
      20'h08391: out <= 12'h660;
      20'h08392: out <= 12'h660;
      20'h08393: out <= 12'h660;
      20'h08394: out <= 12'hbb0;
      20'h08395: out <= 12'h660;
      20'h08396: out <= 12'hee9;
      20'h08397: out <= 12'hee9;
      20'h08398: out <= 12'hbb0;
      20'h08399: out <= 12'hbb0;
      20'h0839a: out <= 12'h660;
      20'h0839b: out <= 12'h660;
      20'h0839c: out <= 12'hbb0;
      20'h0839d: out <= 12'hee9;
      20'h0839e: out <= 12'hbb0;
      20'h0839f: out <= 12'h222;
      20'h083a0: out <= 12'h000;
      20'h083a1: out <= 12'h000;
      20'h083a2: out <= 12'h660;
      20'h083a3: out <= 12'hee9;
      20'h083a4: out <= 12'hbb0;
      20'h083a5: out <= 12'h660;
      20'h083a6: out <= 12'hee9;
      20'h083a7: out <= 12'hee9;
      20'h083a8: out <= 12'hee9;
      20'h083a9: out <= 12'hee9;
      20'h083aa: out <= 12'hee9;
      20'h083ab: out <= 12'h660;
      20'h083ac: out <= 12'hbb0;
      20'h083ad: out <= 12'hee9;
      20'h083ae: out <= 12'h660;
      20'h083af: out <= 12'h000;
      20'h083b0: out <= 12'h222;
      20'h083b1: out <= 12'h222;
      20'h083b2: out <= 12'h660;
      20'h083b3: out <= 12'h660;
      20'h083b4: out <= 12'hbb0;
      20'h083b5: out <= 12'h660;
      20'h083b6: out <= 12'hee9;
      20'h083b7: out <= 12'hee9;
      20'h083b8: out <= 12'hee9;
      20'h083b9: out <= 12'hee9;
      20'h083ba: out <= 12'hee9;
      20'h083bb: out <= 12'h660;
      20'h083bc: out <= 12'hbb0;
      20'h083bd: out <= 12'h660;
      20'h083be: out <= 12'h660;
      20'h083bf: out <= 12'h222;
      20'h083c0: out <= 12'h603;
      20'h083c1: out <= 12'h603;
      20'h083c2: out <= 12'h603;
      20'h083c3: out <= 12'h603;
      20'h083c4: out <= 12'h603;
      20'h083c5: out <= 12'h603;
      20'h083c6: out <= 12'h603;
      20'h083c7: out <= 12'h603;
      20'h083c8: out <= 12'h603;
      20'h083c9: out <= 12'h603;
      20'h083ca: out <= 12'h603;
      20'h083cb: out <= 12'h603;
      20'h083cc: out <= 12'hee9;
      20'h083cd: out <= 12'hee9;
      20'h083ce: out <= 12'hee9;
      20'h083cf: out <= 12'hee9;
      20'h083d0: out <= 12'hee9;
      20'h083d1: out <= 12'hee9;
      20'h083d2: out <= 12'hee9;
      20'h083d3: out <= 12'hb27;
      20'h083d4: out <= 12'hee9;
      20'h083d5: out <= 12'hee9;
      20'h083d6: out <= 12'hee9;
      20'h083d7: out <= 12'hee9;
      20'h083d8: out <= 12'hee9;
      20'h083d9: out <= 12'hee9;
      20'h083da: out <= 12'hee9;
      20'h083db: out <= 12'hb27;
      20'h083dc: out <= 12'hee9;
      20'h083dd: out <= 12'hee9;
      20'h083de: out <= 12'hee9;
      20'h083df: out <= 12'hee9;
      20'h083e0: out <= 12'hee9;
      20'h083e1: out <= 12'hee9;
      20'h083e2: out <= 12'hee9;
      20'h083e3: out <= 12'hb27;
      20'h083e4: out <= 12'hee9;
      20'h083e5: out <= 12'hee9;
      20'h083e6: out <= 12'hee9;
      20'h083e7: out <= 12'hee9;
      20'h083e8: out <= 12'hee9;
      20'h083e9: out <= 12'hee9;
      20'h083ea: out <= 12'hee9;
      20'h083eb: out <= 12'hb27;
      20'h083ec: out <= 12'h603;
      20'h083ed: out <= 12'h603;
      20'h083ee: out <= 12'h603;
      20'h083ef: out <= 12'h603;
      20'h083f0: out <= 12'h603;
      20'h083f1: out <= 12'h603;
      20'h083f2: out <= 12'h603;
      20'h083f3: out <= 12'h603;
      20'h083f4: out <= 12'h603;
      20'h083f5: out <= 12'h603;
      20'h083f6: out <= 12'h603;
      20'h083f7: out <= 12'h603;
      20'h083f8: out <= 12'h603;
      20'h083f9: out <= 12'h603;
      20'h083fa: out <= 12'h603;
      20'h083fb: out <= 12'h603;
      20'h083fc: out <= 12'h603;
      20'h083fd: out <= 12'h603;
      20'h083fe: out <= 12'h603;
      20'h083ff: out <= 12'h603;
      20'h08400: out <= 12'h603;
      20'h08401: out <= 12'h603;
      20'h08402: out <= 12'h603;
      20'h08403: out <= 12'h603;
      20'h08404: out <= 12'h603;
      20'h08405: out <= 12'h603;
      20'h08406: out <= 12'h603;
      20'h08407: out <= 12'h603;
      20'h08408: out <= 12'h603;
      20'h08409: out <= 12'h603;
      20'h0840a: out <= 12'h603;
      20'h0840b: out <= 12'h603;
      20'h0840c: out <= 12'h603;
      20'h0840d: out <= 12'h603;
      20'h0840e: out <= 12'h603;
      20'h0840f: out <= 12'h603;
      20'h08410: out <= 12'h603;
      20'h08411: out <= 12'h603;
      20'h08412: out <= 12'h603;
      20'h08413: out <= 12'h603;
      20'h08414: out <= 12'h603;
      20'h08415: out <= 12'h603;
      20'h08416: out <= 12'h603;
      20'h08417: out <= 12'h603;
      20'h08418: out <= 12'hee9;
      20'h08419: out <= 12'hee9;
      20'h0841a: out <= 12'hee9;
      20'h0841b: out <= 12'hee9;
      20'h0841c: out <= 12'hee9;
      20'h0841d: out <= 12'hee9;
      20'h0841e: out <= 12'hee9;
      20'h0841f: out <= 12'hb27;
      20'h08420: out <= 12'h000;
      20'h08421: out <= 12'h000;
      20'h08422: out <= 12'h000;
      20'h08423: out <= 12'h000;
      20'h08424: out <= 12'h000;
      20'h08425: out <= 12'h000;
      20'h08426: out <= 12'h000;
      20'h08427: out <= 12'h000;
      20'h08428: out <= 12'h000;
      20'h08429: out <= 12'h000;
      20'h0842a: out <= 12'h000;
      20'h0842b: out <= 12'h000;
      20'h0842c: out <= 12'h000;
      20'h0842d: out <= 12'h000;
      20'h0842e: out <= 12'h000;
      20'h0842f: out <= 12'h000;
      20'h08430: out <= 12'h000;
      20'h08431: out <= 12'h000;
      20'h08432: out <= 12'h000;
      20'h08433: out <= 12'h000;
      20'h08434: out <= 12'h000;
      20'h08435: out <= 12'h000;
      20'h08436: out <= 12'h000;
      20'h08437: out <= 12'h000;
      20'h08438: out <= 12'h000;
      20'h08439: out <= 12'h000;
      20'h0843a: out <= 12'h000;
      20'h0843b: out <= 12'h000;
      20'h0843c: out <= 12'h000;
      20'h0843d: out <= 12'h000;
      20'h0843e: out <= 12'h000;
      20'h0843f: out <= 12'h000;
      20'h08440: out <= 12'h000;
      20'h08441: out <= 12'h000;
      20'h08442: out <= 12'h000;
      20'h08443: out <= 12'h000;
      20'h08444: out <= 12'h000;
      20'h08445: out <= 12'h000;
      20'h08446: out <= 12'h000;
      20'h08447: out <= 12'h000;
      20'h08448: out <= 12'h000;
      20'h08449: out <= 12'h000;
      20'h0844a: out <= 12'h000;
      20'h0844b: out <= 12'h000;
      20'h0844c: out <= 12'h000;
      20'h0844d: out <= 12'h000;
      20'h0844e: out <= 12'h000;
      20'h0844f: out <= 12'h000;
      20'h08450: out <= 12'h000;
      20'h08451: out <= 12'h000;
      20'h08452: out <= 12'h000;
      20'h08453: out <= 12'h000;
      20'h08454: out <= 12'h000;
      20'h08455: out <= 12'h000;
      20'h08456: out <= 12'h000;
      20'h08457: out <= 12'h000;
      20'h08458: out <= 12'h000;
      20'h08459: out <= 12'hbb0;
      20'h0845a: out <= 12'hee9;
      20'h0845b: out <= 12'hbb0;
      20'h0845c: out <= 12'h660;
      20'h0845d: out <= 12'h660;
      20'h0845e: out <= 12'hbb0;
      20'h0845f: out <= 12'hbb0;
      20'h08460: out <= 12'hee9;
      20'h08461: out <= 12'hee9;
      20'h08462: out <= 12'h660;
      20'h08463: out <= 12'h660;
      20'h08464: out <= 12'h660;
      20'h08465: out <= 12'hee9;
      20'h08466: out <= 12'hbb0;
      20'h08467: out <= 12'h000;
      20'h08468: out <= 12'h222;
      20'h08469: out <= 12'hbb0;
      20'h0846a: out <= 12'hee9;
      20'h0846b: out <= 12'hbb0;
      20'h0846c: out <= 12'h660;
      20'h0846d: out <= 12'h660;
      20'h0846e: out <= 12'hbb0;
      20'h0846f: out <= 12'hbb0;
      20'h08470: out <= 12'hee9;
      20'h08471: out <= 12'hee9;
      20'h08472: out <= 12'h660;
      20'h08473: out <= 12'h660;
      20'h08474: out <= 12'h660;
      20'h08475: out <= 12'hee9;
      20'h08476: out <= 12'hbb0;
      20'h08477: out <= 12'h222;
      20'h08478: out <= 12'h000;
      20'h08479: out <= 12'h000;
      20'h0847a: out <= 12'h660;
      20'h0847b: out <= 12'hee9;
      20'h0847c: out <= 12'hbb0;
      20'h0847d: out <= 12'h660;
      20'h0847e: out <= 12'hbb0;
      20'h0847f: out <= 12'hbb0;
      20'h08480: out <= 12'hbb0;
      20'h08481: out <= 12'hbb0;
      20'h08482: out <= 12'hbb0;
      20'h08483: out <= 12'h660;
      20'h08484: out <= 12'hbb0;
      20'h08485: out <= 12'hee9;
      20'h08486: out <= 12'h660;
      20'h08487: out <= 12'h000;
      20'h08488: out <= 12'h222;
      20'h08489: out <= 12'h222;
      20'h0848a: out <= 12'h660;
      20'h0848b: out <= 12'h660;
      20'h0848c: out <= 12'hbb0;
      20'h0848d: out <= 12'h660;
      20'h0848e: out <= 12'hbb0;
      20'h0848f: out <= 12'hbb0;
      20'h08490: out <= 12'hbb0;
      20'h08491: out <= 12'hbb0;
      20'h08492: out <= 12'hbb0;
      20'h08493: out <= 12'h660;
      20'h08494: out <= 12'hbb0;
      20'h08495: out <= 12'h660;
      20'h08496: out <= 12'h660;
      20'h08497: out <= 12'h222;
      20'h08498: out <= 12'h000;
      20'h08499: out <= 12'hbb0;
      20'h0849a: out <= 12'hee9;
      20'h0849b: out <= 12'h660;
      20'h0849c: out <= 12'h660;
      20'h0849d: out <= 12'h660;
      20'h0849e: out <= 12'hee9;
      20'h0849f: out <= 12'hee9;
      20'h084a0: out <= 12'hbb0;
      20'h084a1: out <= 12'hbb0;
      20'h084a2: out <= 12'h660;
      20'h084a3: out <= 12'h660;
      20'h084a4: out <= 12'hbb0;
      20'h084a5: out <= 12'hee9;
      20'h084a6: out <= 12'hbb0;
      20'h084a7: out <= 12'h000;
      20'h084a8: out <= 12'h222;
      20'h084a9: out <= 12'hbb0;
      20'h084aa: out <= 12'hee9;
      20'h084ab: out <= 12'h660;
      20'h084ac: out <= 12'h660;
      20'h084ad: out <= 12'h660;
      20'h084ae: out <= 12'hee9;
      20'h084af: out <= 12'hee9;
      20'h084b0: out <= 12'hbb0;
      20'h084b1: out <= 12'hbb0;
      20'h084b2: out <= 12'h660;
      20'h084b3: out <= 12'h660;
      20'h084b4: out <= 12'hbb0;
      20'h084b5: out <= 12'hee9;
      20'h084b6: out <= 12'hbb0;
      20'h084b7: out <= 12'h222;
      20'h084b8: out <= 12'h000;
      20'h084b9: out <= 12'h000;
      20'h084ba: out <= 12'h660;
      20'h084bb: out <= 12'h660;
      20'h084bc: out <= 12'hbb0;
      20'h084bd: out <= 12'h660;
      20'h084be: out <= 12'hee9;
      20'h084bf: out <= 12'hee9;
      20'h084c0: out <= 12'hee9;
      20'h084c1: out <= 12'hee9;
      20'h084c2: out <= 12'hee9;
      20'h084c3: out <= 12'h660;
      20'h084c4: out <= 12'hbb0;
      20'h084c5: out <= 12'h660;
      20'h084c6: out <= 12'h660;
      20'h084c7: out <= 12'h000;
      20'h084c8: out <= 12'h222;
      20'h084c9: out <= 12'h222;
      20'h084ca: out <= 12'h660;
      20'h084cb: out <= 12'hee9;
      20'h084cc: out <= 12'hbb0;
      20'h084cd: out <= 12'h660;
      20'h084ce: out <= 12'hee9;
      20'h084cf: out <= 12'hee9;
      20'h084d0: out <= 12'hee9;
      20'h084d1: out <= 12'hee9;
      20'h084d2: out <= 12'hee9;
      20'h084d3: out <= 12'h660;
      20'h084d4: out <= 12'hbb0;
      20'h084d5: out <= 12'hee9;
      20'h084d6: out <= 12'h660;
      20'h084d7: out <= 12'h222;
      20'h084d8: out <= 12'h603;
      20'h084d9: out <= 12'h603;
      20'h084da: out <= 12'h603;
      20'h084db: out <= 12'h603;
      20'h084dc: out <= 12'h603;
      20'h084dd: out <= 12'h603;
      20'h084de: out <= 12'h603;
      20'h084df: out <= 12'h603;
      20'h084e0: out <= 12'h603;
      20'h084e1: out <= 12'h603;
      20'h084e2: out <= 12'h603;
      20'h084e3: out <= 12'h603;
      20'h084e4: out <= 12'hee9;
      20'h084e5: out <= 12'hf87;
      20'h084e6: out <= 12'hf87;
      20'h084e7: out <= 12'hf87;
      20'h084e8: out <= 12'hf87;
      20'h084e9: out <= 12'hf87;
      20'h084ea: out <= 12'hf87;
      20'h084eb: out <= 12'hb27;
      20'h084ec: out <= 12'hee9;
      20'h084ed: out <= 12'hf87;
      20'h084ee: out <= 12'hf87;
      20'h084ef: out <= 12'hf87;
      20'h084f0: out <= 12'hf87;
      20'h084f1: out <= 12'hf87;
      20'h084f2: out <= 12'hf87;
      20'h084f3: out <= 12'hb27;
      20'h084f4: out <= 12'hee9;
      20'h084f5: out <= 12'hf87;
      20'h084f6: out <= 12'hf87;
      20'h084f7: out <= 12'hf87;
      20'h084f8: out <= 12'hf87;
      20'h084f9: out <= 12'hf87;
      20'h084fa: out <= 12'hf87;
      20'h084fb: out <= 12'hb27;
      20'h084fc: out <= 12'hee9;
      20'h084fd: out <= 12'hf87;
      20'h084fe: out <= 12'hf87;
      20'h084ff: out <= 12'hf87;
      20'h08500: out <= 12'hf87;
      20'h08501: out <= 12'hf87;
      20'h08502: out <= 12'hf87;
      20'h08503: out <= 12'hb27;
      20'h08504: out <= 12'h603;
      20'h08505: out <= 12'h603;
      20'h08506: out <= 12'h603;
      20'h08507: out <= 12'h603;
      20'h08508: out <= 12'h603;
      20'h08509: out <= 12'h603;
      20'h0850a: out <= 12'h603;
      20'h0850b: out <= 12'h603;
      20'h0850c: out <= 12'h603;
      20'h0850d: out <= 12'h603;
      20'h0850e: out <= 12'h603;
      20'h0850f: out <= 12'h603;
      20'h08510: out <= 12'h603;
      20'h08511: out <= 12'h603;
      20'h08512: out <= 12'h603;
      20'h08513: out <= 12'h603;
      20'h08514: out <= 12'h603;
      20'h08515: out <= 12'h603;
      20'h08516: out <= 12'h603;
      20'h08517: out <= 12'h603;
      20'h08518: out <= 12'h603;
      20'h08519: out <= 12'h603;
      20'h0851a: out <= 12'h603;
      20'h0851b: out <= 12'h603;
      20'h0851c: out <= 12'h603;
      20'h0851d: out <= 12'h603;
      20'h0851e: out <= 12'h603;
      20'h0851f: out <= 12'h603;
      20'h08520: out <= 12'h603;
      20'h08521: out <= 12'h603;
      20'h08522: out <= 12'h603;
      20'h08523: out <= 12'h603;
      20'h08524: out <= 12'h603;
      20'h08525: out <= 12'h603;
      20'h08526: out <= 12'h603;
      20'h08527: out <= 12'h603;
      20'h08528: out <= 12'h603;
      20'h08529: out <= 12'h603;
      20'h0852a: out <= 12'h603;
      20'h0852b: out <= 12'h603;
      20'h0852c: out <= 12'h603;
      20'h0852d: out <= 12'h603;
      20'h0852e: out <= 12'h603;
      20'h0852f: out <= 12'h603;
      20'h08530: out <= 12'hee9;
      20'h08531: out <= 12'hf87;
      20'h08532: out <= 12'hf87;
      20'h08533: out <= 12'hf87;
      20'h08534: out <= 12'hf87;
      20'h08535: out <= 12'hf87;
      20'h08536: out <= 12'hf87;
      20'h08537: out <= 12'hb27;
      20'h08538: out <= 12'h000;
      20'h08539: out <= 12'h000;
      20'h0853a: out <= 12'h000;
      20'h0853b: out <= 12'h000;
      20'h0853c: out <= 12'h000;
      20'h0853d: out <= 12'h000;
      20'h0853e: out <= 12'h000;
      20'h0853f: out <= 12'h000;
      20'h08540: out <= 12'h000;
      20'h08541: out <= 12'h000;
      20'h08542: out <= 12'h000;
      20'h08543: out <= 12'h000;
      20'h08544: out <= 12'h000;
      20'h08545: out <= 12'h000;
      20'h08546: out <= 12'h000;
      20'h08547: out <= 12'h000;
      20'h08548: out <= 12'h000;
      20'h08549: out <= 12'h000;
      20'h0854a: out <= 12'h000;
      20'h0854b: out <= 12'h000;
      20'h0854c: out <= 12'h000;
      20'h0854d: out <= 12'h000;
      20'h0854e: out <= 12'h000;
      20'h0854f: out <= 12'h000;
      20'h08550: out <= 12'h000;
      20'h08551: out <= 12'h000;
      20'h08552: out <= 12'h000;
      20'h08553: out <= 12'h000;
      20'h08554: out <= 12'h000;
      20'h08555: out <= 12'h000;
      20'h08556: out <= 12'h000;
      20'h08557: out <= 12'h000;
      20'h08558: out <= 12'h000;
      20'h08559: out <= 12'h000;
      20'h0855a: out <= 12'h000;
      20'h0855b: out <= 12'h000;
      20'h0855c: out <= 12'h000;
      20'h0855d: out <= 12'h000;
      20'h0855e: out <= 12'h000;
      20'h0855f: out <= 12'h000;
      20'h08560: out <= 12'h000;
      20'h08561: out <= 12'h000;
      20'h08562: out <= 12'h000;
      20'h08563: out <= 12'h000;
      20'h08564: out <= 12'h000;
      20'h08565: out <= 12'h000;
      20'h08566: out <= 12'h000;
      20'h08567: out <= 12'h000;
      20'h08568: out <= 12'h000;
      20'h08569: out <= 12'h000;
      20'h0856a: out <= 12'h000;
      20'h0856b: out <= 12'h000;
      20'h0856c: out <= 12'h000;
      20'h0856d: out <= 12'h000;
      20'h0856e: out <= 12'h000;
      20'h0856f: out <= 12'h000;
      20'h08570: out <= 12'h000;
      20'h08571: out <= 12'h660;
      20'h08572: out <= 12'hbb0;
      20'h08573: out <= 12'hee9;
      20'h08574: out <= 12'h660;
      20'h08575: out <= 12'h660;
      20'h08576: out <= 12'h660;
      20'h08577: out <= 12'h660;
      20'h08578: out <= 12'h660;
      20'h08579: out <= 12'h660;
      20'h0857a: out <= 12'hbb0;
      20'h0857b: out <= 12'hbb0;
      20'h0857c: out <= 12'hee9;
      20'h0857d: out <= 12'hbb0;
      20'h0857e: out <= 12'h660;
      20'h0857f: out <= 12'h000;
      20'h08580: out <= 12'h222;
      20'h08581: out <= 12'h660;
      20'h08582: out <= 12'hbb0;
      20'h08583: out <= 12'hee9;
      20'h08584: out <= 12'h660;
      20'h08585: out <= 12'h660;
      20'h08586: out <= 12'h660;
      20'h08587: out <= 12'h660;
      20'h08588: out <= 12'h660;
      20'h08589: out <= 12'h660;
      20'h0858a: out <= 12'h660;
      20'h0858b: out <= 12'hbb0;
      20'h0858c: out <= 12'hee9;
      20'h0858d: out <= 12'hbb0;
      20'h0858e: out <= 12'h660;
      20'h0858f: out <= 12'h222;
      20'h08590: out <= 12'h000;
      20'h08591: out <= 12'h000;
      20'h08592: out <= 12'h660;
      20'h08593: out <= 12'h660;
      20'h08594: out <= 12'hbb0;
      20'h08595: out <= 12'h660;
      20'h08596: out <= 12'h660;
      20'h08597: out <= 12'h660;
      20'h08598: out <= 12'h660;
      20'h08599: out <= 12'h660;
      20'h0859a: out <= 12'h660;
      20'h0859b: out <= 12'h660;
      20'h0859c: out <= 12'hbb0;
      20'h0859d: out <= 12'h660;
      20'h0859e: out <= 12'h660;
      20'h0859f: out <= 12'h000;
      20'h085a0: out <= 12'h222;
      20'h085a1: out <= 12'h222;
      20'h085a2: out <= 12'h660;
      20'h085a3: out <= 12'hee9;
      20'h085a4: out <= 12'hbb0;
      20'h085a5: out <= 12'h660;
      20'h085a6: out <= 12'h660;
      20'h085a7: out <= 12'h660;
      20'h085a8: out <= 12'h660;
      20'h085a9: out <= 12'h660;
      20'h085aa: out <= 12'h660;
      20'h085ab: out <= 12'h660;
      20'h085ac: out <= 12'hbb0;
      20'h085ad: out <= 12'hee9;
      20'h085ae: out <= 12'h660;
      20'h085af: out <= 12'h222;
      20'h085b0: out <= 12'h000;
      20'h085b1: out <= 12'h660;
      20'h085b2: out <= 12'hbb0;
      20'h085b3: out <= 12'hee9;
      20'h085b4: out <= 12'hbb0;
      20'h085b5: out <= 12'hbb0;
      20'h085b6: out <= 12'h660;
      20'h085b7: out <= 12'h660;
      20'h085b8: out <= 12'h660;
      20'h085b9: out <= 12'h660;
      20'h085ba: out <= 12'h660;
      20'h085bb: out <= 12'h660;
      20'h085bc: out <= 12'hee9;
      20'h085bd: out <= 12'hbb0;
      20'h085be: out <= 12'h660;
      20'h085bf: out <= 12'h000;
      20'h085c0: out <= 12'h222;
      20'h085c1: out <= 12'h660;
      20'h085c2: out <= 12'hbb0;
      20'h085c3: out <= 12'hee9;
      20'h085c4: out <= 12'hbb0;
      20'h085c5: out <= 12'h660;
      20'h085c6: out <= 12'h660;
      20'h085c7: out <= 12'h660;
      20'h085c8: out <= 12'h660;
      20'h085c9: out <= 12'h660;
      20'h085ca: out <= 12'h660;
      20'h085cb: out <= 12'h660;
      20'h085cc: out <= 12'hee9;
      20'h085cd: out <= 12'hbb0;
      20'h085ce: out <= 12'h660;
      20'h085cf: out <= 12'h222;
      20'h085d0: out <= 12'h000;
      20'h085d1: out <= 12'h000;
      20'h085d2: out <= 12'h660;
      20'h085d3: out <= 12'hee9;
      20'h085d4: out <= 12'hbb0;
      20'h085d5: out <= 12'hbb0;
      20'h085d6: out <= 12'h660;
      20'h085d7: out <= 12'h660;
      20'h085d8: out <= 12'h660;
      20'h085d9: out <= 12'h660;
      20'h085da: out <= 12'h660;
      20'h085db: out <= 12'hbb0;
      20'h085dc: out <= 12'hbb0;
      20'h085dd: out <= 12'hee9;
      20'h085de: out <= 12'h660;
      20'h085df: out <= 12'h000;
      20'h085e0: out <= 12'h222;
      20'h085e1: out <= 12'h222;
      20'h085e2: out <= 12'h660;
      20'h085e3: out <= 12'h660;
      20'h085e4: out <= 12'hbb0;
      20'h085e5: out <= 12'h660;
      20'h085e6: out <= 12'h660;
      20'h085e7: out <= 12'h660;
      20'h085e8: out <= 12'h660;
      20'h085e9: out <= 12'h660;
      20'h085ea: out <= 12'h660;
      20'h085eb: out <= 12'h660;
      20'h085ec: out <= 12'hbb0;
      20'h085ed: out <= 12'h660;
      20'h085ee: out <= 12'h660;
      20'h085ef: out <= 12'h222;
      20'h085f0: out <= 12'h603;
      20'h085f1: out <= 12'h603;
      20'h085f2: out <= 12'h603;
      20'h085f3: out <= 12'h603;
      20'h085f4: out <= 12'h603;
      20'h085f5: out <= 12'h603;
      20'h085f6: out <= 12'h603;
      20'h085f7: out <= 12'h603;
      20'h085f8: out <= 12'h603;
      20'h085f9: out <= 12'h603;
      20'h085fa: out <= 12'h603;
      20'h085fb: out <= 12'h603;
      20'h085fc: out <= 12'hee9;
      20'h085fd: out <= 12'hf87;
      20'h085fe: out <= 12'hee9;
      20'h085ff: out <= 12'hee9;
      20'h08600: out <= 12'hee9;
      20'h08601: out <= 12'hb27;
      20'h08602: out <= 12'hf87;
      20'h08603: out <= 12'hb27;
      20'h08604: out <= 12'hee9;
      20'h08605: out <= 12'hf87;
      20'h08606: out <= 12'hee9;
      20'h08607: out <= 12'hee9;
      20'h08608: out <= 12'hee9;
      20'h08609: out <= 12'hb27;
      20'h0860a: out <= 12'hf87;
      20'h0860b: out <= 12'hb27;
      20'h0860c: out <= 12'hee9;
      20'h0860d: out <= 12'hf87;
      20'h0860e: out <= 12'hee9;
      20'h0860f: out <= 12'hee9;
      20'h08610: out <= 12'hee9;
      20'h08611: out <= 12'hb27;
      20'h08612: out <= 12'hf87;
      20'h08613: out <= 12'hb27;
      20'h08614: out <= 12'hee9;
      20'h08615: out <= 12'hf87;
      20'h08616: out <= 12'hee9;
      20'h08617: out <= 12'hee9;
      20'h08618: out <= 12'hee9;
      20'h08619: out <= 12'hb27;
      20'h0861a: out <= 12'hf87;
      20'h0861b: out <= 12'hb27;
      20'h0861c: out <= 12'h603;
      20'h0861d: out <= 12'h603;
      20'h0861e: out <= 12'h603;
      20'h0861f: out <= 12'h603;
      20'h08620: out <= 12'h603;
      20'h08621: out <= 12'h603;
      20'h08622: out <= 12'h603;
      20'h08623: out <= 12'h603;
      20'h08624: out <= 12'h603;
      20'h08625: out <= 12'h603;
      20'h08626: out <= 12'h603;
      20'h08627: out <= 12'h603;
      20'h08628: out <= 12'h603;
      20'h08629: out <= 12'h603;
      20'h0862a: out <= 12'h603;
      20'h0862b: out <= 12'h603;
      20'h0862c: out <= 12'h603;
      20'h0862d: out <= 12'h603;
      20'h0862e: out <= 12'h603;
      20'h0862f: out <= 12'h603;
      20'h08630: out <= 12'h603;
      20'h08631: out <= 12'h603;
      20'h08632: out <= 12'h603;
      20'h08633: out <= 12'h603;
      20'h08634: out <= 12'h603;
      20'h08635: out <= 12'h603;
      20'h08636: out <= 12'h603;
      20'h08637: out <= 12'h603;
      20'h08638: out <= 12'h603;
      20'h08639: out <= 12'h603;
      20'h0863a: out <= 12'h603;
      20'h0863b: out <= 12'h603;
      20'h0863c: out <= 12'h603;
      20'h0863d: out <= 12'h603;
      20'h0863e: out <= 12'h603;
      20'h0863f: out <= 12'h603;
      20'h08640: out <= 12'h603;
      20'h08641: out <= 12'h603;
      20'h08642: out <= 12'h603;
      20'h08643: out <= 12'h603;
      20'h08644: out <= 12'h603;
      20'h08645: out <= 12'h603;
      20'h08646: out <= 12'h603;
      20'h08647: out <= 12'h603;
      20'h08648: out <= 12'hee9;
      20'h08649: out <= 12'hf87;
      20'h0864a: out <= 12'hee9;
      20'h0864b: out <= 12'hee9;
      20'h0864c: out <= 12'hee9;
      20'h0864d: out <= 12'hb27;
      20'h0864e: out <= 12'hf87;
      20'h0864f: out <= 12'hb27;
      20'h08650: out <= 12'h000;
      20'h08651: out <= 12'h000;
      20'h08652: out <= 12'h000;
      20'h08653: out <= 12'h000;
      20'h08654: out <= 12'h000;
      20'h08655: out <= 12'h000;
      20'h08656: out <= 12'h000;
      20'h08657: out <= 12'h000;
      20'h08658: out <= 12'h000;
      20'h08659: out <= 12'h000;
      20'h0865a: out <= 12'h000;
      20'h0865b: out <= 12'h000;
      20'h0865c: out <= 12'h000;
      20'h0865d: out <= 12'h000;
      20'h0865e: out <= 12'h000;
      20'h0865f: out <= 12'h000;
      20'h08660: out <= 12'h000;
      20'h08661: out <= 12'h000;
      20'h08662: out <= 12'h000;
      20'h08663: out <= 12'h000;
      20'h08664: out <= 12'h000;
      20'h08665: out <= 12'h000;
      20'h08666: out <= 12'h000;
      20'h08667: out <= 12'h000;
      20'h08668: out <= 12'h000;
      20'h08669: out <= 12'h000;
      20'h0866a: out <= 12'h000;
      20'h0866b: out <= 12'h000;
      20'h0866c: out <= 12'h000;
      20'h0866d: out <= 12'h000;
      20'h0866e: out <= 12'h000;
      20'h0866f: out <= 12'h000;
      20'h08670: out <= 12'h000;
      20'h08671: out <= 12'h000;
      20'h08672: out <= 12'h000;
      20'h08673: out <= 12'h000;
      20'h08674: out <= 12'h000;
      20'h08675: out <= 12'h000;
      20'h08676: out <= 12'h000;
      20'h08677: out <= 12'h000;
      20'h08678: out <= 12'h000;
      20'h08679: out <= 12'h000;
      20'h0867a: out <= 12'h000;
      20'h0867b: out <= 12'h000;
      20'h0867c: out <= 12'h000;
      20'h0867d: out <= 12'h000;
      20'h0867e: out <= 12'h000;
      20'h0867f: out <= 12'h000;
      20'h08680: out <= 12'h000;
      20'h08681: out <= 12'h000;
      20'h08682: out <= 12'h000;
      20'h08683: out <= 12'h000;
      20'h08684: out <= 12'h000;
      20'h08685: out <= 12'h000;
      20'h08686: out <= 12'h000;
      20'h08687: out <= 12'h000;
      20'h08688: out <= 12'h000;
      20'h08689: out <= 12'h000;
      20'h0868a: out <= 12'h660;
      20'h0868b: out <= 12'hbb0;
      20'h0868c: out <= 12'hbb0;
      20'h0868d: out <= 12'hbb0;
      20'h0868e: out <= 12'hbb0;
      20'h0868f: out <= 12'hbb0;
      20'h08690: out <= 12'hbb0;
      20'h08691: out <= 12'hbb0;
      20'h08692: out <= 12'hbb0;
      20'h08693: out <= 12'hbb0;
      20'h08694: out <= 12'hbb0;
      20'h08695: out <= 12'h660;
      20'h08696: out <= 12'h000;
      20'h08697: out <= 12'h000;
      20'h08698: out <= 12'h222;
      20'h08699: out <= 12'h222;
      20'h0869a: out <= 12'h660;
      20'h0869b: out <= 12'hbb0;
      20'h0869c: out <= 12'hbb0;
      20'h0869d: out <= 12'hbb0;
      20'h0869e: out <= 12'hbb0;
      20'h0869f: out <= 12'hbb0;
      20'h086a0: out <= 12'hbb0;
      20'h086a1: out <= 12'hbb0;
      20'h086a2: out <= 12'hbb0;
      20'h086a3: out <= 12'hbb0;
      20'h086a4: out <= 12'hbb0;
      20'h086a5: out <= 12'h660;
      20'h086a6: out <= 12'h222;
      20'h086a7: out <= 12'h222;
      20'h086a8: out <= 12'h000;
      20'h086a9: out <= 12'h000;
      20'h086aa: out <= 12'h660;
      20'h086ab: out <= 12'hee9;
      20'h086ac: out <= 12'hbb0;
      20'h086ad: out <= 12'h660;
      20'h086ae: out <= 12'h660;
      20'h086af: out <= 12'h660;
      20'h086b0: out <= 12'h660;
      20'h086b1: out <= 12'h660;
      20'h086b2: out <= 12'h660;
      20'h086b3: out <= 12'h660;
      20'h086b4: out <= 12'hbb0;
      20'h086b5: out <= 12'hee9;
      20'h086b6: out <= 12'h660;
      20'h086b7: out <= 12'h000;
      20'h086b8: out <= 12'h222;
      20'h086b9: out <= 12'h222;
      20'h086ba: out <= 12'h660;
      20'h086bb: out <= 12'h660;
      20'h086bc: out <= 12'hbb0;
      20'h086bd: out <= 12'h660;
      20'h086be: out <= 12'h660;
      20'h086bf: out <= 12'h660;
      20'h086c0: out <= 12'h660;
      20'h086c1: out <= 12'h660;
      20'h086c2: out <= 12'h660;
      20'h086c3: out <= 12'h660;
      20'h086c4: out <= 12'hbb0;
      20'h086c5: out <= 12'h660;
      20'h086c6: out <= 12'h660;
      20'h086c7: out <= 12'h222;
      20'h086c8: out <= 12'h000;
      20'h086c9: out <= 12'h000;
      20'h086ca: out <= 12'h660;
      20'h086cb: out <= 12'hbb0;
      20'h086cc: out <= 12'hbb0;
      20'h086cd: out <= 12'hbb0;
      20'h086ce: out <= 12'hbb0;
      20'h086cf: out <= 12'hbb0;
      20'h086d0: out <= 12'hbb0;
      20'h086d1: out <= 12'hbb0;
      20'h086d2: out <= 12'hbb0;
      20'h086d3: out <= 12'hbb0;
      20'h086d4: out <= 12'hbb0;
      20'h086d5: out <= 12'h660;
      20'h086d6: out <= 12'h000;
      20'h086d7: out <= 12'h000;
      20'h086d8: out <= 12'h222;
      20'h086d9: out <= 12'h222;
      20'h086da: out <= 12'h660;
      20'h086db: out <= 12'hbb0;
      20'h086dc: out <= 12'hbb0;
      20'h086dd: out <= 12'hbb0;
      20'h086de: out <= 12'hbb0;
      20'h086df: out <= 12'hbb0;
      20'h086e0: out <= 12'hbb0;
      20'h086e1: out <= 12'hbb0;
      20'h086e2: out <= 12'hbb0;
      20'h086e3: out <= 12'hbb0;
      20'h086e4: out <= 12'hbb0;
      20'h086e5: out <= 12'h660;
      20'h086e6: out <= 12'h222;
      20'h086e7: out <= 12'h222;
      20'h086e8: out <= 12'h000;
      20'h086e9: out <= 12'h000;
      20'h086ea: out <= 12'h660;
      20'h086eb: out <= 12'h660;
      20'h086ec: out <= 12'hbb0;
      20'h086ed: out <= 12'hbb0;
      20'h086ee: out <= 12'h660;
      20'h086ef: out <= 12'hbb0;
      20'h086f0: out <= 12'hee9;
      20'h086f1: out <= 12'hbb0;
      20'h086f2: out <= 12'h660;
      20'h086f3: out <= 12'hbb0;
      20'h086f4: out <= 12'hbb0;
      20'h086f5: out <= 12'h660;
      20'h086f6: out <= 12'h660;
      20'h086f7: out <= 12'h000;
      20'h086f8: out <= 12'h222;
      20'h086f9: out <= 12'h222;
      20'h086fa: out <= 12'h660;
      20'h086fb: out <= 12'hee9;
      20'h086fc: out <= 12'hbb0;
      20'h086fd: out <= 12'hbb0;
      20'h086fe: out <= 12'h660;
      20'h086ff: out <= 12'hbb0;
      20'h08700: out <= 12'hee9;
      20'h08701: out <= 12'hbb0;
      20'h08702: out <= 12'h660;
      20'h08703: out <= 12'hbb0;
      20'h08704: out <= 12'hbb0;
      20'h08705: out <= 12'hee9;
      20'h08706: out <= 12'h660;
      20'h08707: out <= 12'h222;
      20'h08708: out <= 12'h603;
      20'h08709: out <= 12'h603;
      20'h0870a: out <= 12'h603;
      20'h0870b: out <= 12'h603;
      20'h0870c: out <= 12'h603;
      20'h0870d: out <= 12'h603;
      20'h0870e: out <= 12'h603;
      20'h0870f: out <= 12'h603;
      20'h08710: out <= 12'h603;
      20'h08711: out <= 12'h603;
      20'h08712: out <= 12'h603;
      20'h08713: out <= 12'h603;
      20'h08714: out <= 12'hee9;
      20'h08715: out <= 12'hf87;
      20'h08716: out <= 12'hee9;
      20'h08717: out <= 12'hf87;
      20'h08718: out <= 12'hf87;
      20'h08719: out <= 12'hb27;
      20'h0871a: out <= 12'hf87;
      20'h0871b: out <= 12'hb27;
      20'h0871c: out <= 12'hee9;
      20'h0871d: out <= 12'hf87;
      20'h0871e: out <= 12'hee9;
      20'h0871f: out <= 12'hf87;
      20'h08720: out <= 12'hf87;
      20'h08721: out <= 12'hb27;
      20'h08722: out <= 12'hf87;
      20'h08723: out <= 12'hb27;
      20'h08724: out <= 12'hee9;
      20'h08725: out <= 12'hf87;
      20'h08726: out <= 12'hee9;
      20'h08727: out <= 12'hf87;
      20'h08728: out <= 12'hf87;
      20'h08729: out <= 12'hb27;
      20'h0872a: out <= 12'hf87;
      20'h0872b: out <= 12'hb27;
      20'h0872c: out <= 12'hee9;
      20'h0872d: out <= 12'hf87;
      20'h0872e: out <= 12'hee9;
      20'h0872f: out <= 12'hf87;
      20'h08730: out <= 12'hf87;
      20'h08731: out <= 12'hb27;
      20'h08732: out <= 12'hf87;
      20'h08733: out <= 12'hb27;
      20'h08734: out <= 12'h603;
      20'h08735: out <= 12'h603;
      20'h08736: out <= 12'h603;
      20'h08737: out <= 12'h603;
      20'h08738: out <= 12'h603;
      20'h08739: out <= 12'h603;
      20'h0873a: out <= 12'h603;
      20'h0873b: out <= 12'h603;
      20'h0873c: out <= 12'h603;
      20'h0873d: out <= 12'h603;
      20'h0873e: out <= 12'h603;
      20'h0873f: out <= 12'h603;
      20'h08740: out <= 12'h603;
      20'h08741: out <= 12'h603;
      20'h08742: out <= 12'h603;
      20'h08743: out <= 12'h603;
      20'h08744: out <= 12'h603;
      20'h08745: out <= 12'h603;
      20'h08746: out <= 12'h603;
      20'h08747: out <= 12'h603;
      20'h08748: out <= 12'h603;
      20'h08749: out <= 12'h603;
      20'h0874a: out <= 12'h603;
      20'h0874b: out <= 12'h603;
      20'h0874c: out <= 12'h603;
      20'h0874d: out <= 12'h603;
      20'h0874e: out <= 12'h603;
      20'h0874f: out <= 12'h603;
      20'h08750: out <= 12'h603;
      20'h08751: out <= 12'h603;
      20'h08752: out <= 12'h603;
      20'h08753: out <= 12'h603;
      20'h08754: out <= 12'h603;
      20'h08755: out <= 12'h603;
      20'h08756: out <= 12'h603;
      20'h08757: out <= 12'h603;
      20'h08758: out <= 12'h603;
      20'h08759: out <= 12'h603;
      20'h0875a: out <= 12'h603;
      20'h0875b: out <= 12'h603;
      20'h0875c: out <= 12'h603;
      20'h0875d: out <= 12'h603;
      20'h0875e: out <= 12'h603;
      20'h0875f: out <= 12'h603;
      20'h08760: out <= 12'hee9;
      20'h08761: out <= 12'hf87;
      20'h08762: out <= 12'hee9;
      20'h08763: out <= 12'hf87;
      20'h08764: out <= 12'hf87;
      20'h08765: out <= 12'hb27;
      20'h08766: out <= 12'hf87;
      20'h08767: out <= 12'hb27;
      20'h08768: out <= 12'h000;
      20'h08769: out <= 12'h000;
      20'h0876a: out <= 12'h000;
      20'h0876b: out <= 12'h000;
      20'h0876c: out <= 12'h000;
      20'h0876d: out <= 12'h000;
      20'h0876e: out <= 12'h000;
      20'h0876f: out <= 12'h000;
      20'h08770: out <= 12'h000;
      20'h08771: out <= 12'h000;
      20'h08772: out <= 12'h000;
      20'h08773: out <= 12'h000;
      20'h08774: out <= 12'h000;
      20'h08775: out <= 12'h000;
      20'h08776: out <= 12'h000;
      20'h08777: out <= 12'h000;
      20'h08778: out <= 12'h000;
      20'h08779: out <= 12'h000;
      20'h0877a: out <= 12'h000;
      20'h0877b: out <= 12'h000;
      20'h0877c: out <= 12'h000;
      20'h0877d: out <= 12'h000;
      20'h0877e: out <= 12'h000;
      20'h0877f: out <= 12'h000;
      20'h08780: out <= 12'h000;
      20'h08781: out <= 12'h000;
      20'h08782: out <= 12'h000;
      20'h08783: out <= 12'h000;
      20'h08784: out <= 12'h000;
      20'h08785: out <= 12'h000;
      20'h08786: out <= 12'h000;
      20'h08787: out <= 12'h000;
      20'h08788: out <= 12'h000;
      20'h08789: out <= 12'h000;
      20'h0878a: out <= 12'h000;
      20'h0878b: out <= 12'h000;
      20'h0878c: out <= 12'h000;
      20'h0878d: out <= 12'h000;
      20'h0878e: out <= 12'h000;
      20'h0878f: out <= 12'h000;
      20'h08790: out <= 12'h000;
      20'h08791: out <= 12'h000;
      20'h08792: out <= 12'h000;
      20'h08793: out <= 12'h000;
      20'h08794: out <= 12'h000;
      20'h08795: out <= 12'h000;
      20'h08796: out <= 12'h000;
      20'h08797: out <= 12'h000;
      20'h08798: out <= 12'h000;
      20'h08799: out <= 12'h000;
      20'h0879a: out <= 12'h000;
      20'h0879b: out <= 12'h000;
      20'h0879c: out <= 12'h000;
      20'h0879d: out <= 12'h000;
      20'h0879e: out <= 12'h000;
      20'h0879f: out <= 12'h000;
      20'h087a0: out <= 12'h000;
      20'h087a1: out <= 12'h000;
      20'h087a2: out <= 12'hee9;
      20'h087a3: out <= 12'h660;
      20'h087a4: out <= 12'hee9;
      20'h087a5: out <= 12'h660;
      20'h087a6: out <= 12'hee9;
      20'h087a7: out <= 12'h660;
      20'h087a8: out <= 12'hee9;
      20'h087a9: out <= 12'h660;
      20'h087aa: out <= 12'hee9;
      20'h087ab: out <= 12'h660;
      20'h087ac: out <= 12'hee9;
      20'h087ad: out <= 12'h660;
      20'h087ae: out <= 12'h000;
      20'h087af: out <= 12'h000;
      20'h087b0: out <= 12'h222;
      20'h087b1: out <= 12'h222;
      20'h087b2: out <= 12'h660;
      20'h087b3: out <= 12'hee9;
      20'h087b4: out <= 12'h660;
      20'h087b5: out <= 12'hee9;
      20'h087b6: out <= 12'h660;
      20'h087b7: out <= 12'hee9;
      20'h087b8: out <= 12'h660;
      20'h087b9: out <= 12'hee9;
      20'h087ba: out <= 12'h660;
      20'h087bb: out <= 12'hee9;
      20'h087bc: out <= 12'h660;
      20'h087bd: out <= 12'hee9;
      20'h087be: out <= 12'h222;
      20'h087bf: out <= 12'h222;
      20'h087c0: out <= 12'h000;
      20'h087c1: out <= 12'h000;
      20'h087c2: out <= 12'h660;
      20'h087c3: out <= 12'h660;
      20'h087c4: out <= 12'hbb0;
      20'h087c5: out <= 12'hee9;
      20'h087c6: out <= 12'hbb0;
      20'h087c7: out <= 12'hbb0;
      20'h087c8: out <= 12'hbb0;
      20'h087c9: out <= 12'hbb0;
      20'h087ca: out <= 12'hbb0;
      20'h087cb: out <= 12'hee9;
      20'h087cc: out <= 12'hbb0;
      20'h087cd: out <= 12'h660;
      20'h087ce: out <= 12'h660;
      20'h087cf: out <= 12'h000;
      20'h087d0: out <= 12'h222;
      20'h087d1: out <= 12'h222;
      20'h087d2: out <= 12'h660;
      20'h087d3: out <= 12'hee9;
      20'h087d4: out <= 12'hbb0;
      20'h087d5: out <= 12'hee9;
      20'h087d6: out <= 12'hbb0;
      20'h087d7: out <= 12'hbb0;
      20'h087d8: out <= 12'hbb0;
      20'h087d9: out <= 12'hbb0;
      20'h087da: out <= 12'hbb0;
      20'h087db: out <= 12'hee9;
      20'h087dc: out <= 12'hbb0;
      20'h087dd: out <= 12'hee9;
      20'h087de: out <= 12'h660;
      20'h087df: out <= 12'h222;
      20'h087e0: out <= 12'h000;
      20'h087e1: out <= 12'h000;
      20'h087e2: out <= 12'h660;
      20'h087e3: out <= 12'hee9;
      20'h087e4: out <= 12'h660;
      20'h087e5: out <= 12'hee9;
      20'h087e6: out <= 12'h660;
      20'h087e7: out <= 12'hee9;
      20'h087e8: out <= 12'h660;
      20'h087e9: out <= 12'hee9;
      20'h087ea: out <= 12'h660;
      20'h087eb: out <= 12'hee9;
      20'h087ec: out <= 12'h660;
      20'h087ed: out <= 12'hee9;
      20'h087ee: out <= 12'h000;
      20'h087ef: out <= 12'h000;
      20'h087f0: out <= 12'h222;
      20'h087f1: out <= 12'h222;
      20'h087f2: out <= 12'hee9;
      20'h087f3: out <= 12'h660;
      20'h087f4: out <= 12'hee9;
      20'h087f5: out <= 12'h660;
      20'h087f6: out <= 12'hee9;
      20'h087f7: out <= 12'h660;
      20'h087f8: out <= 12'hee9;
      20'h087f9: out <= 12'h660;
      20'h087fa: out <= 12'hee9;
      20'h087fb: out <= 12'h660;
      20'h087fc: out <= 12'hee9;
      20'h087fd: out <= 12'h660;
      20'h087fe: out <= 12'h222;
      20'h087ff: out <= 12'h222;
      20'h08800: out <= 12'h000;
      20'h08801: out <= 12'h000;
      20'h08802: out <= 12'h660;
      20'h08803: out <= 12'hee9;
      20'h08804: out <= 12'hbb0;
      20'h08805: out <= 12'hee9;
      20'h08806: out <= 12'h660;
      20'h08807: out <= 12'h660;
      20'h08808: out <= 12'hee9;
      20'h08809: out <= 12'h660;
      20'h0880a: out <= 12'h660;
      20'h0880b: out <= 12'hee9;
      20'h0880c: out <= 12'hbb0;
      20'h0880d: out <= 12'hee9;
      20'h0880e: out <= 12'h660;
      20'h0880f: out <= 12'h000;
      20'h08810: out <= 12'h222;
      20'h08811: out <= 12'h222;
      20'h08812: out <= 12'h660;
      20'h08813: out <= 12'h660;
      20'h08814: out <= 12'hbb0;
      20'h08815: out <= 12'hee9;
      20'h08816: out <= 12'h660;
      20'h08817: out <= 12'h660;
      20'h08818: out <= 12'hee9;
      20'h08819: out <= 12'h660;
      20'h0881a: out <= 12'h660;
      20'h0881b: out <= 12'hee9;
      20'h0881c: out <= 12'hbb0;
      20'h0881d: out <= 12'h660;
      20'h0881e: out <= 12'h660;
      20'h0881f: out <= 12'h222;
      20'h08820: out <= 12'h603;
      20'h08821: out <= 12'h603;
      20'h08822: out <= 12'h603;
      20'h08823: out <= 12'h603;
      20'h08824: out <= 12'h603;
      20'h08825: out <= 12'h603;
      20'h08826: out <= 12'h603;
      20'h08827: out <= 12'h603;
      20'h08828: out <= 12'h603;
      20'h08829: out <= 12'h603;
      20'h0882a: out <= 12'h603;
      20'h0882b: out <= 12'h603;
      20'h0882c: out <= 12'hee9;
      20'h0882d: out <= 12'hf87;
      20'h0882e: out <= 12'hee9;
      20'h0882f: out <= 12'hf87;
      20'h08830: out <= 12'hf87;
      20'h08831: out <= 12'hb27;
      20'h08832: out <= 12'hf87;
      20'h08833: out <= 12'hb27;
      20'h08834: out <= 12'hee9;
      20'h08835: out <= 12'hf87;
      20'h08836: out <= 12'hee9;
      20'h08837: out <= 12'hf87;
      20'h08838: out <= 12'hf87;
      20'h08839: out <= 12'hb27;
      20'h0883a: out <= 12'hf87;
      20'h0883b: out <= 12'hb27;
      20'h0883c: out <= 12'hee9;
      20'h0883d: out <= 12'hf87;
      20'h0883e: out <= 12'hee9;
      20'h0883f: out <= 12'hf87;
      20'h08840: out <= 12'hf87;
      20'h08841: out <= 12'hb27;
      20'h08842: out <= 12'hf87;
      20'h08843: out <= 12'hb27;
      20'h08844: out <= 12'hee9;
      20'h08845: out <= 12'hf87;
      20'h08846: out <= 12'hee9;
      20'h08847: out <= 12'hf87;
      20'h08848: out <= 12'hf87;
      20'h08849: out <= 12'hb27;
      20'h0884a: out <= 12'hf87;
      20'h0884b: out <= 12'hb27;
      20'h0884c: out <= 12'h603;
      20'h0884d: out <= 12'h603;
      20'h0884e: out <= 12'h603;
      20'h0884f: out <= 12'h603;
      20'h08850: out <= 12'h603;
      20'h08851: out <= 12'h603;
      20'h08852: out <= 12'h603;
      20'h08853: out <= 12'h603;
      20'h08854: out <= 12'h603;
      20'h08855: out <= 12'h603;
      20'h08856: out <= 12'h603;
      20'h08857: out <= 12'h603;
      20'h08858: out <= 12'h603;
      20'h08859: out <= 12'h603;
      20'h0885a: out <= 12'h603;
      20'h0885b: out <= 12'h603;
      20'h0885c: out <= 12'h603;
      20'h0885d: out <= 12'h603;
      20'h0885e: out <= 12'h603;
      20'h0885f: out <= 12'h603;
      20'h08860: out <= 12'h603;
      20'h08861: out <= 12'h603;
      20'h08862: out <= 12'h603;
      20'h08863: out <= 12'h603;
      20'h08864: out <= 12'h603;
      20'h08865: out <= 12'h603;
      20'h08866: out <= 12'h603;
      20'h08867: out <= 12'h603;
      20'h08868: out <= 12'h603;
      20'h08869: out <= 12'h603;
      20'h0886a: out <= 12'h603;
      20'h0886b: out <= 12'h603;
      20'h0886c: out <= 12'h603;
      20'h0886d: out <= 12'h603;
      20'h0886e: out <= 12'h603;
      20'h0886f: out <= 12'h603;
      20'h08870: out <= 12'h603;
      20'h08871: out <= 12'h603;
      20'h08872: out <= 12'h603;
      20'h08873: out <= 12'h603;
      20'h08874: out <= 12'h603;
      20'h08875: out <= 12'h603;
      20'h08876: out <= 12'h603;
      20'h08877: out <= 12'h603;
      20'h08878: out <= 12'hee9;
      20'h08879: out <= 12'hf87;
      20'h0887a: out <= 12'hee9;
      20'h0887b: out <= 12'hf87;
      20'h0887c: out <= 12'hf87;
      20'h0887d: out <= 12'hb27;
      20'h0887e: out <= 12'hf87;
      20'h0887f: out <= 12'hb27;
      20'h08880: out <= 12'h000;
      20'h08881: out <= 12'h000;
      20'h08882: out <= 12'h000;
      20'h08883: out <= 12'h000;
      20'h08884: out <= 12'h000;
      20'h08885: out <= 12'h000;
      20'h08886: out <= 12'h000;
      20'h08887: out <= 12'h000;
      20'h08888: out <= 12'h000;
      20'h08889: out <= 12'h000;
      20'h0888a: out <= 12'h000;
      20'h0888b: out <= 12'h000;
      20'h0888c: out <= 12'h000;
      20'h0888d: out <= 12'h000;
      20'h0888e: out <= 12'h000;
      20'h0888f: out <= 12'h000;
      20'h08890: out <= 12'h000;
      20'h08891: out <= 12'h000;
      20'h08892: out <= 12'h000;
      20'h08893: out <= 12'h000;
      20'h08894: out <= 12'h000;
      20'h08895: out <= 12'h000;
      20'h08896: out <= 12'h000;
      20'h08897: out <= 12'h000;
      20'h08898: out <= 12'h000;
      20'h08899: out <= 12'h000;
      20'h0889a: out <= 12'h000;
      20'h0889b: out <= 12'h000;
      20'h0889c: out <= 12'h000;
      20'h0889d: out <= 12'h000;
      20'h0889e: out <= 12'h000;
      20'h0889f: out <= 12'h000;
      20'h088a0: out <= 12'h000;
      20'h088a1: out <= 12'h000;
      20'h088a2: out <= 12'h000;
      20'h088a3: out <= 12'h000;
      20'h088a4: out <= 12'h000;
      20'h088a5: out <= 12'h000;
      20'h088a6: out <= 12'h000;
      20'h088a7: out <= 12'h000;
      20'h088a8: out <= 12'h000;
      20'h088a9: out <= 12'h000;
      20'h088aa: out <= 12'h000;
      20'h088ab: out <= 12'h000;
      20'h088ac: out <= 12'h000;
      20'h088ad: out <= 12'h000;
      20'h088ae: out <= 12'h000;
      20'h088af: out <= 12'h000;
      20'h088b0: out <= 12'h000;
      20'h088b1: out <= 12'h000;
      20'h088b2: out <= 12'h000;
      20'h088b3: out <= 12'h000;
      20'h088b4: out <= 12'h000;
      20'h088b5: out <= 12'h000;
      20'h088b6: out <= 12'h000;
      20'h088b7: out <= 12'h000;
      20'h088b8: out <= 12'h000;
      20'h088b9: out <= 12'h000;
      20'h088ba: out <= 12'h660;
      20'h088bb: out <= 12'h660;
      20'h088bc: out <= 12'h660;
      20'h088bd: out <= 12'h660;
      20'h088be: out <= 12'h660;
      20'h088bf: out <= 12'h660;
      20'h088c0: out <= 12'h660;
      20'h088c1: out <= 12'h660;
      20'h088c2: out <= 12'h660;
      20'h088c3: out <= 12'h660;
      20'h088c4: out <= 12'h660;
      20'h088c5: out <= 12'h660;
      20'h088c6: out <= 12'h000;
      20'h088c7: out <= 12'h000;
      20'h088c8: out <= 12'h222;
      20'h088c9: out <= 12'h222;
      20'h088ca: out <= 12'h660;
      20'h088cb: out <= 12'h660;
      20'h088cc: out <= 12'h660;
      20'h088cd: out <= 12'h660;
      20'h088ce: out <= 12'h660;
      20'h088cf: out <= 12'h660;
      20'h088d0: out <= 12'h660;
      20'h088d1: out <= 12'h660;
      20'h088d2: out <= 12'h660;
      20'h088d3: out <= 12'h660;
      20'h088d4: out <= 12'h660;
      20'h088d5: out <= 12'h660;
      20'h088d6: out <= 12'h222;
      20'h088d7: out <= 12'h222;
      20'h088d8: out <= 12'h000;
      20'h088d9: out <= 12'h000;
      20'h088da: out <= 12'h660;
      20'h088db: out <= 12'hee9;
      20'h088dc: out <= 12'h660;
      20'h088dd: out <= 12'hbb0;
      20'h088de: out <= 12'hee9;
      20'h088df: out <= 12'hee9;
      20'h088e0: out <= 12'hee9;
      20'h088e1: out <= 12'hee9;
      20'h088e2: out <= 12'hee9;
      20'h088e3: out <= 12'hbb0;
      20'h088e4: out <= 12'h660;
      20'h088e5: out <= 12'hee9;
      20'h088e6: out <= 12'h660;
      20'h088e7: out <= 12'h000;
      20'h088e8: out <= 12'h222;
      20'h088e9: out <= 12'h222;
      20'h088ea: out <= 12'h660;
      20'h088eb: out <= 12'h660;
      20'h088ec: out <= 12'h660;
      20'h088ed: out <= 12'hbb0;
      20'h088ee: out <= 12'hee9;
      20'h088ef: out <= 12'hee9;
      20'h088f0: out <= 12'hee9;
      20'h088f1: out <= 12'hee9;
      20'h088f2: out <= 12'hee9;
      20'h088f3: out <= 12'hbb0;
      20'h088f4: out <= 12'h660;
      20'h088f5: out <= 12'h660;
      20'h088f6: out <= 12'h660;
      20'h088f7: out <= 12'h222;
      20'h088f8: out <= 12'h000;
      20'h088f9: out <= 12'h000;
      20'h088fa: out <= 12'h660;
      20'h088fb: out <= 12'h660;
      20'h088fc: out <= 12'h660;
      20'h088fd: out <= 12'h660;
      20'h088fe: out <= 12'h660;
      20'h088ff: out <= 12'h660;
      20'h08900: out <= 12'h660;
      20'h08901: out <= 12'h660;
      20'h08902: out <= 12'h660;
      20'h08903: out <= 12'h660;
      20'h08904: out <= 12'h660;
      20'h08905: out <= 12'h660;
      20'h08906: out <= 12'h000;
      20'h08907: out <= 12'h000;
      20'h08908: out <= 12'h222;
      20'h08909: out <= 12'h222;
      20'h0890a: out <= 12'h660;
      20'h0890b: out <= 12'h660;
      20'h0890c: out <= 12'h660;
      20'h0890d: out <= 12'h660;
      20'h0890e: out <= 12'h660;
      20'h0890f: out <= 12'h660;
      20'h08910: out <= 12'h660;
      20'h08911: out <= 12'h660;
      20'h08912: out <= 12'h660;
      20'h08913: out <= 12'h660;
      20'h08914: out <= 12'h660;
      20'h08915: out <= 12'h660;
      20'h08916: out <= 12'h222;
      20'h08917: out <= 12'h222;
      20'h08918: out <= 12'h000;
      20'h08919: out <= 12'h000;
      20'h0891a: out <= 12'h660;
      20'h0891b: out <= 12'h660;
      20'h0891c: out <= 12'h660;
      20'h0891d: out <= 12'hbb0;
      20'h0891e: out <= 12'hee9;
      20'h0891f: out <= 12'h660;
      20'h08920: out <= 12'hee9;
      20'h08921: out <= 12'h660;
      20'h08922: out <= 12'hee9;
      20'h08923: out <= 12'hbb0;
      20'h08924: out <= 12'h660;
      20'h08925: out <= 12'h660;
      20'h08926: out <= 12'h660;
      20'h08927: out <= 12'h000;
      20'h08928: out <= 12'h222;
      20'h08929: out <= 12'h222;
      20'h0892a: out <= 12'h660;
      20'h0892b: out <= 12'hee9;
      20'h0892c: out <= 12'h660;
      20'h0892d: out <= 12'hbb0;
      20'h0892e: out <= 12'hee9;
      20'h0892f: out <= 12'h660;
      20'h08930: out <= 12'hee9;
      20'h08931: out <= 12'h660;
      20'h08932: out <= 12'hee9;
      20'h08933: out <= 12'hbb0;
      20'h08934: out <= 12'h660;
      20'h08935: out <= 12'hee9;
      20'h08936: out <= 12'h660;
      20'h08937: out <= 12'h222;
      20'h08938: out <= 12'h603;
      20'h08939: out <= 12'h603;
      20'h0893a: out <= 12'h603;
      20'h0893b: out <= 12'h603;
      20'h0893c: out <= 12'h603;
      20'h0893d: out <= 12'h603;
      20'h0893e: out <= 12'h603;
      20'h0893f: out <= 12'h603;
      20'h08940: out <= 12'h603;
      20'h08941: out <= 12'h603;
      20'h08942: out <= 12'h603;
      20'h08943: out <= 12'h603;
      20'h08944: out <= 12'hee9;
      20'h08945: out <= 12'hf87;
      20'h08946: out <= 12'hee9;
      20'h08947: out <= 12'hb27;
      20'h08948: out <= 12'hb27;
      20'h08949: out <= 12'hb27;
      20'h0894a: out <= 12'hf87;
      20'h0894b: out <= 12'hb27;
      20'h0894c: out <= 12'hee9;
      20'h0894d: out <= 12'hf87;
      20'h0894e: out <= 12'hee9;
      20'h0894f: out <= 12'hb27;
      20'h08950: out <= 12'hb27;
      20'h08951: out <= 12'hb27;
      20'h08952: out <= 12'hf87;
      20'h08953: out <= 12'hb27;
      20'h08954: out <= 12'hee9;
      20'h08955: out <= 12'hf87;
      20'h08956: out <= 12'hee9;
      20'h08957: out <= 12'hb27;
      20'h08958: out <= 12'hb27;
      20'h08959: out <= 12'hb27;
      20'h0895a: out <= 12'hf87;
      20'h0895b: out <= 12'hb27;
      20'h0895c: out <= 12'hee9;
      20'h0895d: out <= 12'hf87;
      20'h0895e: out <= 12'hee9;
      20'h0895f: out <= 12'hb27;
      20'h08960: out <= 12'hb27;
      20'h08961: out <= 12'hb27;
      20'h08962: out <= 12'hf87;
      20'h08963: out <= 12'hb27;
      20'h08964: out <= 12'h603;
      20'h08965: out <= 12'h603;
      20'h08966: out <= 12'h603;
      20'h08967: out <= 12'h603;
      20'h08968: out <= 12'h603;
      20'h08969: out <= 12'h603;
      20'h0896a: out <= 12'h603;
      20'h0896b: out <= 12'h603;
      20'h0896c: out <= 12'h603;
      20'h0896d: out <= 12'h603;
      20'h0896e: out <= 12'h603;
      20'h0896f: out <= 12'h603;
      20'h08970: out <= 12'h603;
      20'h08971: out <= 12'h603;
      20'h08972: out <= 12'h603;
      20'h08973: out <= 12'h603;
      20'h08974: out <= 12'h603;
      20'h08975: out <= 12'h603;
      20'h08976: out <= 12'h603;
      20'h08977: out <= 12'h603;
      20'h08978: out <= 12'h603;
      20'h08979: out <= 12'h603;
      20'h0897a: out <= 12'h603;
      20'h0897b: out <= 12'h603;
      20'h0897c: out <= 12'h603;
      20'h0897d: out <= 12'h603;
      20'h0897e: out <= 12'h603;
      20'h0897f: out <= 12'h603;
      20'h08980: out <= 12'h603;
      20'h08981: out <= 12'h603;
      20'h08982: out <= 12'h603;
      20'h08983: out <= 12'h603;
      20'h08984: out <= 12'h603;
      20'h08985: out <= 12'h603;
      20'h08986: out <= 12'h603;
      20'h08987: out <= 12'h603;
      20'h08988: out <= 12'h603;
      20'h08989: out <= 12'h603;
      20'h0898a: out <= 12'h603;
      20'h0898b: out <= 12'h603;
      20'h0898c: out <= 12'h603;
      20'h0898d: out <= 12'h603;
      20'h0898e: out <= 12'h603;
      20'h0898f: out <= 12'h603;
      20'h08990: out <= 12'hee9;
      20'h08991: out <= 12'hf87;
      20'h08992: out <= 12'hee9;
      20'h08993: out <= 12'hb27;
      20'h08994: out <= 12'hb27;
      20'h08995: out <= 12'hb27;
      20'h08996: out <= 12'hf87;
      20'h08997: out <= 12'hb27;
      20'h08998: out <= 12'h000;
      20'h08999: out <= 12'h000;
      20'h0899a: out <= 12'h000;
      20'h0899b: out <= 12'h000;
      20'h0899c: out <= 12'h000;
      20'h0899d: out <= 12'h000;
      20'h0899e: out <= 12'h000;
      20'h0899f: out <= 12'h000;
      20'h089a0: out <= 12'h000;
      20'h089a1: out <= 12'h000;
      20'h089a2: out <= 12'h000;
      20'h089a3: out <= 12'h000;
      20'h089a4: out <= 12'h000;
      20'h089a5: out <= 12'h000;
      20'h089a6: out <= 12'h000;
      20'h089a7: out <= 12'h000;
      20'h089a8: out <= 12'h000;
      20'h089a9: out <= 12'h000;
      20'h089aa: out <= 12'h000;
      20'h089ab: out <= 12'h000;
      20'h089ac: out <= 12'h000;
      20'h089ad: out <= 12'h000;
      20'h089ae: out <= 12'h000;
      20'h089af: out <= 12'h000;
      20'h089b0: out <= 12'h000;
      20'h089b1: out <= 12'h000;
      20'h089b2: out <= 12'h000;
      20'h089b3: out <= 12'h000;
      20'h089b4: out <= 12'h000;
      20'h089b5: out <= 12'h000;
      20'h089b6: out <= 12'h000;
      20'h089b7: out <= 12'h000;
      20'h089b8: out <= 12'h000;
      20'h089b9: out <= 12'h000;
      20'h089ba: out <= 12'h000;
      20'h089bb: out <= 12'h000;
      20'h089bc: out <= 12'h000;
      20'h089bd: out <= 12'h000;
      20'h089be: out <= 12'h000;
      20'h089bf: out <= 12'h000;
      20'h089c0: out <= 12'h000;
      20'h089c1: out <= 12'h000;
      20'h089c2: out <= 12'h000;
      20'h089c3: out <= 12'h000;
      20'h089c4: out <= 12'h000;
      20'h089c5: out <= 12'h000;
      20'h089c6: out <= 12'h000;
      20'h089c7: out <= 12'h000;
      20'h089c8: out <= 12'h000;
      20'h089c9: out <= 12'h000;
      20'h089ca: out <= 12'h000;
      20'h089cb: out <= 12'h000;
      20'h089cc: out <= 12'h000;
      20'h089cd: out <= 12'h000;
      20'h089ce: out <= 12'h000;
      20'h089cf: out <= 12'h000;
      20'h089d0: out <= 12'h000;
      20'h089d1: out <= 12'h000;
      20'h089d2: out <= 12'h000;
      20'h089d3: out <= 12'h000;
      20'h089d4: out <= 12'h000;
      20'h089d5: out <= 12'h000;
      20'h089d6: out <= 12'h000;
      20'h089d7: out <= 12'h000;
      20'h089d8: out <= 12'h000;
      20'h089d9: out <= 12'h000;
      20'h089da: out <= 12'h000;
      20'h089db: out <= 12'h000;
      20'h089dc: out <= 12'h000;
      20'h089dd: out <= 12'h000;
      20'h089de: out <= 12'h000;
      20'h089df: out <= 12'h000;
      20'h089e0: out <= 12'h222;
      20'h089e1: out <= 12'h222;
      20'h089e2: out <= 12'h222;
      20'h089e3: out <= 12'h222;
      20'h089e4: out <= 12'h222;
      20'h089e5: out <= 12'h222;
      20'h089e6: out <= 12'h222;
      20'h089e7: out <= 12'h222;
      20'h089e8: out <= 12'h222;
      20'h089e9: out <= 12'h222;
      20'h089ea: out <= 12'h222;
      20'h089eb: out <= 12'h222;
      20'h089ec: out <= 12'h222;
      20'h089ed: out <= 12'h222;
      20'h089ee: out <= 12'h222;
      20'h089ef: out <= 12'h222;
      20'h089f0: out <= 12'h000;
      20'h089f1: out <= 12'h000;
      20'h089f2: out <= 12'h000;
      20'h089f3: out <= 12'h000;
      20'h089f4: out <= 12'h000;
      20'h089f5: out <= 12'h660;
      20'h089f6: out <= 12'hbb0;
      20'h089f7: out <= 12'hbb0;
      20'h089f8: out <= 12'hbb0;
      20'h089f9: out <= 12'hbb0;
      20'h089fa: out <= 12'hbb0;
      20'h089fb: out <= 12'h660;
      20'h089fc: out <= 12'h000;
      20'h089fd: out <= 12'h000;
      20'h089fe: out <= 12'h000;
      20'h089ff: out <= 12'h000;
      20'h08a00: out <= 12'h222;
      20'h08a01: out <= 12'h222;
      20'h08a02: out <= 12'h222;
      20'h08a03: out <= 12'h222;
      20'h08a04: out <= 12'h222;
      20'h08a05: out <= 12'h660;
      20'h08a06: out <= 12'hbb0;
      20'h08a07: out <= 12'hbb0;
      20'h08a08: out <= 12'hbb0;
      20'h08a09: out <= 12'hbb0;
      20'h08a0a: out <= 12'hbb0;
      20'h08a0b: out <= 12'h660;
      20'h08a0c: out <= 12'h222;
      20'h08a0d: out <= 12'h222;
      20'h08a0e: out <= 12'h222;
      20'h08a0f: out <= 12'h222;
      20'h08a10: out <= 12'h000;
      20'h08a11: out <= 12'h000;
      20'h08a12: out <= 12'h000;
      20'h08a13: out <= 12'h000;
      20'h08a14: out <= 12'h000;
      20'h08a15: out <= 12'h000;
      20'h08a16: out <= 12'h000;
      20'h08a17: out <= 12'h000;
      20'h08a18: out <= 12'h000;
      20'h08a19: out <= 12'h000;
      20'h08a1a: out <= 12'h000;
      20'h08a1b: out <= 12'h000;
      20'h08a1c: out <= 12'h000;
      20'h08a1d: out <= 12'h000;
      20'h08a1e: out <= 12'h000;
      20'h08a1f: out <= 12'h000;
      20'h08a20: out <= 12'h222;
      20'h08a21: out <= 12'h222;
      20'h08a22: out <= 12'h222;
      20'h08a23: out <= 12'h222;
      20'h08a24: out <= 12'h222;
      20'h08a25: out <= 12'h222;
      20'h08a26: out <= 12'h222;
      20'h08a27: out <= 12'h222;
      20'h08a28: out <= 12'h222;
      20'h08a29: out <= 12'h222;
      20'h08a2a: out <= 12'h222;
      20'h08a2b: out <= 12'h222;
      20'h08a2c: out <= 12'h222;
      20'h08a2d: out <= 12'h222;
      20'h08a2e: out <= 12'h222;
      20'h08a2f: out <= 12'h222;
      20'h08a30: out <= 12'h000;
      20'h08a31: out <= 12'h000;
      20'h08a32: out <= 12'h000;
      20'h08a33: out <= 12'h000;
      20'h08a34: out <= 12'h000;
      20'h08a35: out <= 12'h660;
      20'h08a36: out <= 12'hbb0;
      20'h08a37: out <= 12'h660;
      20'h08a38: out <= 12'hee9;
      20'h08a39: out <= 12'h660;
      20'h08a3a: out <= 12'hbb0;
      20'h08a3b: out <= 12'h660;
      20'h08a3c: out <= 12'h000;
      20'h08a3d: out <= 12'h000;
      20'h08a3e: out <= 12'h000;
      20'h08a3f: out <= 12'h000;
      20'h08a40: out <= 12'h222;
      20'h08a41: out <= 12'h222;
      20'h08a42: out <= 12'h222;
      20'h08a43: out <= 12'h222;
      20'h08a44: out <= 12'h222;
      20'h08a45: out <= 12'h660;
      20'h08a46: out <= 12'hbb0;
      20'h08a47: out <= 12'h660;
      20'h08a48: out <= 12'hee9;
      20'h08a49: out <= 12'h660;
      20'h08a4a: out <= 12'hbb0;
      20'h08a4b: out <= 12'h660;
      20'h08a4c: out <= 12'h222;
      20'h08a4d: out <= 12'h222;
      20'h08a4e: out <= 12'h222;
      20'h08a4f: out <= 12'h222;
      20'h08a50: out <= 12'h603;
      20'h08a51: out <= 12'h603;
      20'h08a52: out <= 12'h603;
      20'h08a53: out <= 12'h603;
      20'h08a54: out <= 12'h603;
      20'h08a55: out <= 12'h603;
      20'h08a56: out <= 12'h603;
      20'h08a57: out <= 12'h603;
      20'h08a58: out <= 12'h603;
      20'h08a59: out <= 12'h603;
      20'h08a5a: out <= 12'h603;
      20'h08a5b: out <= 12'h603;
      20'h08a5c: out <= 12'hee9;
      20'h08a5d: out <= 12'hf87;
      20'h08a5e: out <= 12'hf87;
      20'h08a5f: out <= 12'hf87;
      20'h08a60: out <= 12'hf87;
      20'h08a61: out <= 12'hf87;
      20'h08a62: out <= 12'hf87;
      20'h08a63: out <= 12'hb27;
      20'h08a64: out <= 12'hee9;
      20'h08a65: out <= 12'hf87;
      20'h08a66: out <= 12'hf87;
      20'h08a67: out <= 12'hf87;
      20'h08a68: out <= 12'hf87;
      20'h08a69: out <= 12'hf87;
      20'h08a6a: out <= 12'hf87;
      20'h08a6b: out <= 12'hb27;
      20'h08a6c: out <= 12'hee9;
      20'h08a6d: out <= 12'hf87;
      20'h08a6e: out <= 12'hf87;
      20'h08a6f: out <= 12'hf87;
      20'h08a70: out <= 12'hf87;
      20'h08a71: out <= 12'hf87;
      20'h08a72: out <= 12'hf87;
      20'h08a73: out <= 12'hb27;
      20'h08a74: out <= 12'hee9;
      20'h08a75: out <= 12'hf87;
      20'h08a76: out <= 12'hf87;
      20'h08a77: out <= 12'hf87;
      20'h08a78: out <= 12'hf87;
      20'h08a79: out <= 12'hf87;
      20'h08a7a: out <= 12'hf87;
      20'h08a7b: out <= 12'hb27;
      20'h08a7c: out <= 12'h603;
      20'h08a7d: out <= 12'h603;
      20'h08a7e: out <= 12'h603;
      20'h08a7f: out <= 12'h603;
      20'h08a80: out <= 12'h603;
      20'h08a81: out <= 12'h603;
      20'h08a82: out <= 12'h603;
      20'h08a83: out <= 12'h603;
      20'h08a84: out <= 12'h603;
      20'h08a85: out <= 12'h603;
      20'h08a86: out <= 12'h603;
      20'h08a87: out <= 12'h603;
      20'h08a88: out <= 12'h603;
      20'h08a89: out <= 12'h603;
      20'h08a8a: out <= 12'h603;
      20'h08a8b: out <= 12'h603;
      20'h08a8c: out <= 12'h603;
      20'h08a8d: out <= 12'h603;
      20'h08a8e: out <= 12'h603;
      20'h08a8f: out <= 12'h603;
      20'h08a90: out <= 12'h603;
      20'h08a91: out <= 12'h603;
      20'h08a92: out <= 12'h603;
      20'h08a93: out <= 12'h603;
      20'h08a94: out <= 12'h603;
      20'h08a95: out <= 12'h603;
      20'h08a96: out <= 12'h603;
      20'h08a97: out <= 12'h603;
      20'h08a98: out <= 12'h603;
      20'h08a99: out <= 12'h603;
      20'h08a9a: out <= 12'h603;
      20'h08a9b: out <= 12'h603;
      20'h08a9c: out <= 12'h603;
      20'h08a9d: out <= 12'h603;
      20'h08a9e: out <= 12'h603;
      20'h08a9f: out <= 12'h603;
      20'h08aa0: out <= 12'h603;
      20'h08aa1: out <= 12'h603;
      20'h08aa2: out <= 12'h603;
      20'h08aa3: out <= 12'h603;
      20'h08aa4: out <= 12'h603;
      20'h08aa5: out <= 12'h603;
      20'h08aa6: out <= 12'h603;
      20'h08aa7: out <= 12'h603;
      20'h08aa8: out <= 12'hee9;
      20'h08aa9: out <= 12'hf87;
      20'h08aaa: out <= 12'hf87;
      20'h08aab: out <= 12'hf87;
      20'h08aac: out <= 12'hf87;
      20'h08aad: out <= 12'hf87;
      20'h08aae: out <= 12'hf87;
      20'h08aaf: out <= 12'hb27;
      20'h08ab0: out <= 12'h000;
      20'h08ab1: out <= 12'h000;
      20'h08ab2: out <= 12'h000;
      20'h08ab3: out <= 12'h000;
      20'h08ab4: out <= 12'h000;
      20'h08ab5: out <= 12'h000;
      20'h08ab6: out <= 12'h000;
      20'h08ab7: out <= 12'h000;
      20'h08ab8: out <= 12'h000;
      20'h08ab9: out <= 12'h000;
      20'h08aba: out <= 12'h000;
      20'h08abb: out <= 12'h000;
      20'h08abc: out <= 12'h000;
      20'h08abd: out <= 12'h000;
      20'h08abe: out <= 12'h000;
      20'h08abf: out <= 12'h000;
      20'h08ac0: out <= 12'h000;
      20'h08ac1: out <= 12'h000;
      20'h08ac2: out <= 12'h000;
      20'h08ac3: out <= 12'h000;
      20'h08ac4: out <= 12'h000;
      20'h08ac5: out <= 12'h000;
      20'h08ac6: out <= 12'h000;
      20'h08ac7: out <= 12'h000;
      20'h08ac8: out <= 12'h000;
      20'h08ac9: out <= 12'h000;
      20'h08aca: out <= 12'h000;
      20'h08acb: out <= 12'h000;
      20'h08acc: out <= 12'h000;
      20'h08acd: out <= 12'h000;
      20'h08ace: out <= 12'h000;
      20'h08acf: out <= 12'h000;
      20'h08ad0: out <= 12'h000;
      20'h08ad1: out <= 12'h000;
      20'h08ad2: out <= 12'h000;
      20'h08ad3: out <= 12'h000;
      20'h08ad4: out <= 12'h000;
      20'h08ad5: out <= 12'h000;
      20'h08ad6: out <= 12'h000;
      20'h08ad7: out <= 12'h000;
      20'h08ad8: out <= 12'h000;
      20'h08ad9: out <= 12'h000;
      20'h08ada: out <= 12'h000;
      20'h08adb: out <= 12'h000;
      20'h08adc: out <= 12'h000;
      20'h08add: out <= 12'h000;
      20'h08ade: out <= 12'h000;
      20'h08adf: out <= 12'h000;
      20'h08ae0: out <= 12'h000;
      20'h08ae1: out <= 12'h000;
      20'h08ae2: out <= 12'h000;
      20'h08ae3: out <= 12'h000;
      20'h08ae4: out <= 12'h000;
      20'h08ae5: out <= 12'h000;
      20'h08ae6: out <= 12'h000;
      20'h08ae7: out <= 12'h000;
      20'h08ae8: out <= 12'h000;
      20'h08ae9: out <= 12'h000;
      20'h08aea: out <= 12'h000;
      20'h08aeb: out <= 12'h000;
      20'h08aec: out <= 12'h000;
      20'h08aed: out <= 12'h000;
      20'h08aee: out <= 12'h000;
      20'h08aef: out <= 12'h000;
      20'h08af0: out <= 12'h000;
      20'h08af1: out <= 12'h000;
      20'h08af2: out <= 12'h000;
      20'h08af3: out <= 12'h000;
      20'h08af4: out <= 12'h000;
      20'h08af5: out <= 12'h000;
      20'h08af6: out <= 12'h000;
      20'h08af7: out <= 12'h000;
      20'h08af8: out <= 12'h222;
      20'h08af9: out <= 12'h222;
      20'h08afa: out <= 12'h222;
      20'h08afb: out <= 12'h222;
      20'h08afc: out <= 12'h222;
      20'h08afd: out <= 12'h222;
      20'h08afe: out <= 12'h222;
      20'h08aff: out <= 12'h222;
      20'h08b00: out <= 12'h222;
      20'h08b01: out <= 12'h222;
      20'h08b02: out <= 12'h222;
      20'h08b03: out <= 12'h222;
      20'h08b04: out <= 12'h222;
      20'h08b05: out <= 12'h222;
      20'h08b06: out <= 12'h222;
      20'h08b07: out <= 12'h222;
      20'h08b08: out <= 12'h000;
      20'h08b09: out <= 12'h000;
      20'h08b0a: out <= 12'h000;
      20'h08b0b: out <= 12'h000;
      20'h08b0c: out <= 12'h000;
      20'h08b0d: out <= 12'h000;
      20'h08b0e: out <= 12'h000;
      20'h08b0f: out <= 12'h000;
      20'h08b10: out <= 12'h000;
      20'h08b11: out <= 12'h000;
      20'h08b12: out <= 12'h000;
      20'h08b13: out <= 12'h000;
      20'h08b14: out <= 12'h000;
      20'h08b15: out <= 12'h000;
      20'h08b16: out <= 12'h000;
      20'h08b17: out <= 12'h000;
      20'h08b18: out <= 12'h222;
      20'h08b19: out <= 12'h222;
      20'h08b1a: out <= 12'h222;
      20'h08b1b: out <= 12'h222;
      20'h08b1c: out <= 12'h222;
      20'h08b1d: out <= 12'h222;
      20'h08b1e: out <= 12'h222;
      20'h08b1f: out <= 12'h222;
      20'h08b20: out <= 12'h222;
      20'h08b21: out <= 12'h222;
      20'h08b22: out <= 12'h222;
      20'h08b23: out <= 12'h222;
      20'h08b24: out <= 12'h222;
      20'h08b25: out <= 12'h222;
      20'h08b26: out <= 12'h222;
      20'h08b27: out <= 12'h222;
      20'h08b28: out <= 12'h000;
      20'h08b29: out <= 12'h000;
      20'h08b2a: out <= 12'h000;
      20'h08b2b: out <= 12'h000;
      20'h08b2c: out <= 12'h000;
      20'h08b2d: out <= 12'h000;
      20'h08b2e: out <= 12'h000;
      20'h08b2f: out <= 12'h000;
      20'h08b30: out <= 12'h000;
      20'h08b31: out <= 12'h000;
      20'h08b32: out <= 12'h000;
      20'h08b33: out <= 12'h000;
      20'h08b34: out <= 12'h000;
      20'h08b35: out <= 12'h000;
      20'h08b36: out <= 12'h000;
      20'h08b37: out <= 12'h000;
      20'h08b38: out <= 12'h222;
      20'h08b39: out <= 12'h222;
      20'h08b3a: out <= 12'h222;
      20'h08b3b: out <= 12'h222;
      20'h08b3c: out <= 12'h222;
      20'h08b3d: out <= 12'h222;
      20'h08b3e: out <= 12'h222;
      20'h08b3f: out <= 12'h222;
      20'h08b40: out <= 12'h222;
      20'h08b41: out <= 12'h222;
      20'h08b42: out <= 12'h222;
      20'h08b43: out <= 12'h222;
      20'h08b44: out <= 12'h222;
      20'h08b45: out <= 12'h222;
      20'h08b46: out <= 12'h222;
      20'h08b47: out <= 12'h222;
      20'h08b48: out <= 12'h000;
      20'h08b49: out <= 12'h000;
      20'h08b4a: out <= 12'h000;
      20'h08b4b: out <= 12'h000;
      20'h08b4c: out <= 12'h000;
      20'h08b4d: out <= 12'h000;
      20'h08b4e: out <= 12'h000;
      20'h08b4f: out <= 12'h660;
      20'h08b50: out <= 12'hee9;
      20'h08b51: out <= 12'h660;
      20'h08b52: out <= 12'h000;
      20'h08b53: out <= 12'h000;
      20'h08b54: out <= 12'h000;
      20'h08b55: out <= 12'h000;
      20'h08b56: out <= 12'h000;
      20'h08b57: out <= 12'h000;
      20'h08b58: out <= 12'h222;
      20'h08b59: out <= 12'h222;
      20'h08b5a: out <= 12'h222;
      20'h08b5b: out <= 12'h222;
      20'h08b5c: out <= 12'h222;
      20'h08b5d: out <= 12'h222;
      20'h08b5e: out <= 12'h222;
      20'h08b5f: out <= 12'h660;
      20'h08b60: out <= 12'hee9;
      20'h08b61: out <= 12'h660;
      20'h08b62: out <= 12'h222;
      20'h08b63: out <= 12'h222;
      20'h08b64: out <= 12'h222;
      20'h08b65: out <= 12'h222;
      20'h08b66: out <= 12'h222;
      20'h08b67: out <= 12'h222;
      20'h08b68: out <= 12'h603;
      20'h08b69: out <= 12'h603;
      20'h08b6a: out <= 12'h603;
      20'h08b6b: out <= 12'h603;
      20'h08b6c: out <= 12'h603;
      20'h08b6d: out <= 12'h603;
      20'h08b6e: out <= 12'h603;
      20'h08b6f: out <= 12'h603;
      20'h08b70: out <= 12'h603;
      20'h08b71: out <= 12'h603;
      20'h08b72: out <= 12'h603;
      20'h08b73: out <= 12'h603;
      20'h08b74: out <= 12'hb27;
      20'h08b75: out <= 12'hb27;
      20'h08b76: out <= 12'hb27;
      20'h08b77: out <= 12'hb27;
      20'h08b78: out <= 12'hb27;
      20'h08b79: out <= 12'hb27;
      20'h08b7a: out <= 12'hb27;
      20'h08b7b: out <= 12'hb27;
      20'h08b7c: out <= 12'hb27;
      20'h08b7d: out <= 12'hb27;
      20'h08b7e: out <= 12'hb27;
      20'h08b7f: out <= 12'hb27;
      20'h08b80: out <= 12'hb27;
      20'h08b81: out <= 12'hb27;
      20'h08b82: out <= 12'hb27;
      20'h08b83: out <= 12'hb27;
      20'h08b84: out <= 12'hb27;
      20'h08b85: out <= 12'hb27;
      20'h08b86: out <= 12'hb27;
      20'h08b87: out <= 12'hb27;
      20'h08b88: out <= 12'hb27;
      20'h08b89: out <= 12'hb27;
      20'h08b8a: out <= 12'hb27;
      20'h08b8b: out <= 12'hb27;
      20'h08b8c: out <= 12'hb27;
      20'h08b8d: out <= 12'hb27;
      20'h08b8e: out <= 12'hb27;
      20'h08b8f: out <= 12'hb27;
      20'h08b90: out <= 12'hb27;
      20'h08b91: out <= 12'hb27;
      20'h08b92: out <= 12'hb27;
      20'h08b93: out <= 12'hb27;
      20'h08b94: out <= 12'h603;
      20'h08b95: out <= 12'h603;
      20'h08b96: out <= 12'h603;
      20'h08b97: out <= 12'h603;
      20'h08b98: out <= 12'h603;
      20'h08b99: out <= 12'h603;
      20'h08b9a: out <= 12'h603;
      20'h08b9b: out <= 12'h603;
      20'h08b9c: out <= 12'h603;
      20'h08b9d: out <= 12'h603;
      20'h08b9e: out <= 12'h603;
      20'h08b9f: out <= 12'h603;
      20'h08ba0: out <= 12'h603;
      20'h08ba1: out <= 12'h603;
      20'h08ba2: out <= 12'h603;
      20'h08ba3: out <= 12'h603;
      20'h08ba4: out <= 12'h603;
      20'h08ba5: out <= 12'h603;
      20'h08ba6: out <= 12'h603;
      20'h08ba7: out <= 12'h603;
      20'h08ba8: out <= 12'h603;
      20'h08ba9: out <= 12'h603;
      20'h08baa: out <= 12'h603;
      20'h08bab: out <= 12'h603;
      20'h08bac: out <= 12'h603;
      20'h08bad: out <= 12'h603;
      20'h08bae: out <= 12'h603;
      20'h08baf: out <= 12'h603;
      20'h08bb0: out <= 12'h603;
      20'h08bb1: out <= 12'h603;
      20'h08bb2: out <= 12'h603;
      20'h08bb3: out <= 12'h603;
      20'h08bb4: out <= 12'h603;
      20'h08bb5: out <= 12'h603;
      20'h08bb6: out <= 12'h603;
      20'h08bb7: out <= 12'h603;
      20'h08bb8: out <= 12'h603;
      20'h08bb9: out <= 12'h603;
      20'h08bba: out <= 12'h603;
      20'h08bbb: out <= 12'h603;
      20'h08bbc: out <= 12'h603;
      20'h08bbd: out <= 12'h603;
      20'h08bbe: out <= 12'h603;
      20'h08bbf: out <= 12'h603;
      20'h08bc0: out <= 12'hb27;
      20'h08bc1: out <= 12'hb27;
      20'h08bc2: out <= 12'hb27;
      20'h08bc3: out <= 12'hb27;
      20'h08bc4: out <= 12'hb27;
      20'h08bc5: out <= 12'hb27;
      20'h08bc6: out <= 12'hb27;
      20'h08bc7: out <= 12'hb27;
      20'h08bc8: out <= 12'h000;
      20'h08bc9: out <= 12'h000;
      20'h08bca: out <= 12'h000;
      20'h08bcb: out <= 12'h000;
      20'h08bcc: out <= 12'h000;
      20'h08bcd: out <= 12'h000;
      20'h08bce: out <= 12'h000;
      20'h08bcf: out <= 12'h000;
      20'h08bd0: out <= 12'h000;
      20'h08bd1: out <= 12'h000;
      20'h08bd2: out <= 12'h000;
      20'h08bd3: out <= 12'h000;
      20'h08bd4: out <= 12'h000;
      20'h08bd5: out <= 12'h000;
      20'h08bd6: out <= 12'h000;
      20'h08bd7: out <= 12'h000;
      20'h08bd8: out <= 12'h000;
      20'h08bd9: out <= 12'h000;
      20'h08bda: out <= 12'h000;
      20'h08bdb: out <= 12'h000;
      20'h08bdc: out <= 12'h000;
      20'h08bdd: out <= 12'h000;
      20'h08bde: out <= 12'h000;
      20'h08bdf: out <= 12'h000;
      20'h08be0: out <= 12'h000;
      20'h08be1: out <= 12'h000;
      20'h08be2: out <= 12'h000;
      20'h08be3: out <= 12'h000;
      20'h08be4: out <= 12'h000;
      20'h08be5: out <= 12'h000;
      20'h08be6: out <= 12'h000;
      20'h08be7: out <= 12'h000;
      20'h08be8: out <= 12'h000;
      20'h08be9: out <= 12'h000;
      20'h08bea: out <= 12'h000;
      20'h08beb: out <= 12'h000;
      20'h08bec: out <= 12'h000;
      20'h08bed: out <= 12'h000;
      20'h08bee: out <= 12'h000;
      20'h08bef: out <= 12'h000;
      20'h08bf0: out <= 12'h000;
      20'h08bf1: out <= 12'h000;
      20'h08bf2: out <= 12'h000;
      20'h08bf3: out <= 12'h000;
      20'h08bf4: out <= 12'h000;
      20'h08bf5: out <= 12'h000;
      20'h08bf6: out <= 12'h000;
      20'h08bf7: out <= 12'h000;
      20'h08bf8: out <= 12'h000;
      20'h08bf9: out <= 12'h000;
      20'h08bfa: out <= 12'h000;
      20'h08bfb: out <= 12'h000;
      20'h08bfc: out <= 12'h000;
      20'h08bfd: out <= 12'h000;
      20'h08bfe: out <= 12'h000;
      20'h08bff: out <= 12'h000;
      20'h08c00: out <= 12'h222;
      20'h08c01: out <= 12'h666;
      20'h08c02: out <= 12'h666;
      20'h08c03: out <= 12'h666;
      20'h08c04: out <= 12'h666;
      20'h08c05: out <= 12'h666;
      20'h08c06: out <= 12'h666;
      20'h08c07: out <= 12'h666;
      20'h08c08: out <= 12'h666;
      20'h08c09: out <= 12'h666;
      20'h08c0a: out <= 12'h666;
      20'h08c0b: out <= 12'h666;
      20'h08c0c: out <= 12'h666;
      20'h08c0d: out <= 12'h666;
      20'h08c0e: out <= 12'h666;
      20'h08c0f: out <= 12'h222;
      20'h08c10: out <= 12'h000;
      20'h08c11: out <= 12'h666;
      20'h08c12: out <= 12'h666;
      20'h08c13: out <= 12'h666;
      20'h08c14: out <= 12'h666;
      20'h08c15: out <= 12'h666;
      20'h08c16: out <= 12'h666;
      20'h08c17: out <= 12'h666;
      20'h08c18: out <= 12'h666;
      20'h08c19: out <= 12'h666;
      20'h08c1a: out <= 12'h666;
      20'h08c1b: out <= 12'h666;
      20'h08c1c: out <= 12'h666;
      20'h08c1d: out <= 12'h666;
      20'h08c1e: out <= 12'h666;
      20'h08c1f: out <= 12'h000;
      20'h08c20: out <= 12'h222;
      20'h08c21: out <= 12'h222;
      20'h08c22: out <= 12'h222;
      20'h08c23: out <= 12'h222;
      20'h08c24: out <= 12'h222;
      20'h08c25: out <= 12'h222;
      20'h08c26: out <= 12'hbbb;
      20'h08c27: out <= 12'hbbb;
      20'h08c28: out <= 12'hfff;
      20'h08c29: out <= 12'hbbb;
      20'h08c2a: out <= 12'hbbb;
      20'h08c2b: out <= 12'h222;
      20'h08c2c: out <= 12'h222;
      20'h08c2d: out <= 12'h222;
      20'h08c2e: out <= 12'h222;
      20'h08c2f: out <= 12'h222;
      20'h08c30: out <= 12'h000;
      20'h08c31: out <= 12'h000;
      20'h08c32: out <= 12'h000;
      20'h08c33: out <= 12'h000;
      20'h08c34: out <= 12'h000;
      20'h08c35: out <= 12'h000;
      20'h08c36: out <= 12'hbbb;
      20'h08c37: out <= 12'hbbb;
      20'h08c38: out <= 12'hfff;
      20'h08c39: out <= 12'hbbb;
      20'h08c3a: out <= 12'hbbb;
      20'h08c3b: out <= 12'h000;
      20'h08c3c: out <= 12'h000;
      20'h08c3d: out <= 12'h000;
      20'h08c3e: out <= 12'h000;
      20'h08c3f: out <= 12'h000;
      20'h08c40: out <= 12'h222;
      20'h08c41: out <= 12'h666;
      20'h08c42: out <= 12'h666;
      20'h08c43: out <= 12'h666;
      20'h08c44: out <= 12'h666;
      20'h08c45: out <= 12'h666;
      20'h08c46: out <= 12'h666;
      20'h08c47: out <= 12'h666;
      20'h08c48: out <= 12'h666;
      20'h08c49: out <= 12'h666;
      20'h08c4a: out <= 12'h666;
      20'h08c4b: out <= 12'h666;
      20'h08c4c: out <= 12'h666;
      20'h08c4d: out <= 12'h666;
      20'h08c4e: out <= 12'h666;
      20'h08c4f: out <= 12'h222;
      20'h08c50: out <= 12'h000;
      20'h08c51: out <= 12'h666;
      20'h08c52: out <= 12'h666;
      20'h08c53: out <= 12'h666;
      20'h08c54: out <= 12'h666;
      20'h08c55: out <= 12'h666;
      20'h08c56: out <= 12'h666;
      20'h08c57: out <= 12'h666;
      20'h08c58: out <= 12'h666;
      20'h08c59: out <= 12'h666;
      20'h08c5a: out <= 12'h666;
      20'h08c5b: out <= 12'h666;
      20'h08c5c: out <= 12'h666;
      20'h08c5d: out <= 12'h666;
      20'h08c5e: out <= 12'h666;
      20'h08c5f: out <= 12'h000;
      20'h08c60: out <= 12'h222;
      20'h08c61: out <= 12'h222;
      20'h08c62: out <= 12'h222;
      20'h08c63: out <= 12'h222;
      20'h08c64: out <= 12'h222;
      20'h08c65: out <= 12'h222;
      20'h08c66: out <= 12'h222;
      20'h08c67: out <= 12'h222;
      20'h08c68: out <= 12'h222;
      20'h08c69: out <= 12'h222;
      20'h08c6a: out <= 12'h222;
      20'h08c6b: out <= 12'h222;
      20'h08c6c: out <= 12'h222;
      20'h08c6d: out <= 12'h222;
      20'h08c6e: out <= 12'h222;
      20'h08c6f: out <= 12'h222;
      20'h08c70: out <= 12'h000;
      20'h08c71: out <= 12'h000;
      20'h08c72: out <= 12'h000;
      20'h08c73: out <= 12'h000;
      20'h08c74: out <= 12'h000;
      20'h08c75: out <= 12'h000;
      20'h08c76: out <= 12'h000;
      20'h08c77: out <= 12'h000;
      20'h08c78: out <= 12'h000;
      20'h08c79: out <= 12'h000;
      20'h08c7a: out <= 12'h000;
      20'h08c7b: out <= 12'h000;
      20'h08c7c: out <= 12'h000;
      20'h08c7d: out <= 12'h000;
      20'h08c7e: out <= 12'h000;
      20'h08c7f: out <= 12'h000;
      20'h08c80: out <= 12'h603;
      20'h08c81: out <= 12'h603;
      20'h08c82: out <= 12'h603;
      20'h08c83: out <= 12'h603;
      20'h08c84: out <= 12'h603;
      20'h08c85: out <= 12'h603;
      20'h08c86: out <= 12'h603;
      20'h08c87: out <= 12'h603;
      20'h08c88: out <= 12'h603;
      20'h08c89: out <= 12'h603;
      20'h08c8a: out <= 12'h603;
      20'h08c8b: out <= 12'h603;
      20'h08c8c: out <= 12'h603;
      20'h08c8d: out <= 12'h603;
      20'h08c8e: out <= 12'h603;
      20'h08c8f: out <= 12'h603;
      20'h08c90: out <= 12'h603;
      20'h08c91: out <= 12'h603;
      20'h08c92: out <= 12'h603;
      20'h08c93: out <= 12'h603;
      20'h08c94: out <= 12'h603;
      20'h08c95: out <= 12'h603;
      20'h08c96: out <= 12'h603;
      20'h08c97: out <= 12'h603;
      20'h08c98: out <= 12'h603;
      20'h08c99: out <= 12'h603;
      20'h08c9a: out <= 12'h603;
      20'h08c9b: out <= 12'h603;
      20'h08c9c: out <= 12'h603;
      20'h08c9d: out <= 12'h603;
      20'h08c9e: out <= 12'h603;
      20'h08c9f: out <= 12'h603;
      20'h08ca0: out <= 12'h603;
      20'h08ca1: out <= 12'h603;
      20'h08ca2: out <= 12'h603;
      20'h08ca3: out <= 12'h603;
      20'h08ca4: out <= 12'h603;
      20'h08ca5: out <= 12'h603;
      20'h08ca6: out <= 12'h603;
      20'h08ca7: out <= 12'h603;
      20'h08ca8: out <= 12'h603;
      20'h08ca9: out <= 12'h603;
      20'h08caa: out <= 12'h603;
      20'h08cab: out <= 12'h603;
      20'h08cac: out <= 12'h603;
      20'h08cad: out <= 12'h603;
      20'h08cae: out <= 12'h603;
      20'h08caf: out <= 12'h603;
      20'h08cb0: out <= 12'h603;
      20'h08cb1: out <= 12'h603;
      20'h08cb2: out <= 12'h603;
      20'h08cb3: out <= 12'h603;
      20'h08cb4: out <= 12'h603;
      20'h08cb5: out <= 12'h603;
      20'h08cb6: out <= 12'h603;
      20'h08cb7: out <= 12'h603;
      20'h08cb8: out <= 12'h603;
      20'h08cb9: out <= 12'h603;
      20'h08cba: out <= 12'h603;
      20'h08cbb: out <= 12'h603;
      20'h08cbc: out <= 12'h603;
      20'h08cbd: out <= 12'h603;
      20'h08cbe: out <= 12'h603;
      20'h08cbf: out <= 12'h603;
      20'h08cc0: out <= 12'h603;
      20'h08cc1: out <= 12'h603;
      20'h08cc2: out <= 12'h603;
      20'h08cc3: out <= 12'h603;
      20'h08cc4: out <= 12'h603;
      20'h08cc5: out <= 12'h603;
      20'h08cc6: out <= 12'h603;
      20'h08cc7: out <= 12'h603;
      20'h08cc8: out <= 12'h603;
      20'h08cc9: out <= 12'h603;
      20'h08cca: out <= 12'h603;
      20'h08ccb: out <= 12'h603;
      20'h08ccc: out <= 12'h603;
      20'h08ccd: out <= 12'h603;
      20'h08cce: out <= 12'h603;
      20'h08ccf: out <= 12'h603;
      20'h08cd0: out <= 12'h603;
      20'h08cd1: out <= 12'h603;
      20'h08cd2: out <= 12'h603;
      20'h08cd3: out <= 12'h603;
      20'h08cd4: out <= 12'h603;
      20'h08cd5: out <= 12'h603;
      20'h08cd6: out <= 12'h603;
      20'h08cd7: out <= 12'h603;
      20'h08cd8: out <= 12'hee9;
      20'h08cd9: out <= 12'hee9;
      20'h08cda: out <= 12'hee9;
      20'h08cdb: out <= 12'hee9;
      20'h08cdc: out <= 12'hee9;
      20'h08cdd: out <= 12'hee9;
      20'h08cde: out <= 12'hee9;
      20'h08cdf: out <= 12'hb27;
      20'h08ce0: out <= 12'h000;
      20'h08ce1: out <= 12'h000;
      20'h08ce2: out <= 12'h000;
      20'h08ce3: out <= 12'h000;
      20'h08ce4: out <= 12'h000;
      20'h08ce5: out <= 12'h000;
      20'h08ce6: out <= 12'h000;
      20'h08ce7: out <= 12'h000;
      20'h08ce8: out <= 12'h000;
      20'h08ce9: out <= 12'h8d0;
      20'h08cea: out <= 12'h8d0;
      20'h08ceb: out <= 12'h8d0;
      20'h08cec: out <= 12'h8d0;
      20'h08ced: out <= 12'h8d0;
      20'h08cee: out <= 12'h000;
      20'h08cef: out <= 12'h000;
      20'h08cf0: out <= 12'h8d0;
      20'h08cf1: out <= 12'h8d0;
      20'h08cf2: out <= 12'h8d0;
      20'h08cf3: out <= 12'h8d0;
      20'h08cf4: out <= 12'h8d0;
      20'h08cf5: out <= 12'h000;
      20'h08cf6: out <= 12'h000;
      20'h08cf7: out <= 12'h8d0;
      20'h08cf8: out <= 12'h8d0;
      20'h08cf9: out <= 12'h000;
      20'h08cfa: out <= 12'h000;
      20'h08cfb: out <= 12'h000;
      20'h08cfc: out <= 12'h000;
      20'h08cfd: out <= 12'h000;
      20'h08cfe: out <= 12'h8d0;
      20'h08cff: out <= 12'h8d0;
      20'h08d00: out <= 12'h8d0;
      20'h08d01: out <= 12'h8d0;
      20'h08d02: out <= 12'h000;
      20'h08d03: out <= 12'h000;
      20'h08d04: out <= 12'h8d0;
      20'h08d05: out <= 12'h8d0;
      20'h08d06: out <= 12'h000;
      20'h08d07: out <= 12'h000;
      20'h08d08: out <= 12'h000;
      20'h08d09: out <= 12'h8d0;
      20'h08d0a: out <= 12'h8d0;
      20'h08d0b: out <= 12'h000;
      20'h08d0c: out <= 12'h000;
      20'h08d0d: out <= 12'h000;
      20'h08d0e: out <= 12'h000;
      20'h08d0f: out <= 12'h000;
      20'h08d10: out <= 12'h000;
      20'h08d11: out <= 12'h000;
      20'h08d12: out <= 12'h000;
      20'h08d13: out <= 12'h000;
      20'h08d14: out <= 12'h000;
      20'h08d15: out <= 12'h000;
      20'h08d16: out <= 12'h000;
      20'h08d17: out <= 12'h000;
      20'h08d18: out <= 12'h222;
      20'h08d19: out <= 12'hfff;
      20'h08d1a: out <= 12'h666;
      20'h08d1b: out <= 12'hfff;
      20'h08d1c: out <= 12'h666;
      20'h08d1d: out <= 12'hfff;
      20'h08d1e: out <= 12'h666;
      20'h08d1f: out <= 12'hfff;
      20'h08d20: out <= 12'h666;
      20'h08d21: out <= 12'hfff;
      20'h08d22: out <= 12'h666;
      20'h08d23: out <= 12'hfff;
      20'h08d24: out <= 12'h666;
      20'h08d25: out <= 12'hfff;
      20'h08d26: out <= 12'h666;
      20'h08d27: out <= 12'h222;
      20'h08d28: out <= 12'h000;
      20'h08d29: out <= 12'h666;
      20'h08d2a: out <= 12'hfff;
      20'h08d2b: out <= 12'h666;
      20'h08d2c: out <= 12'hfff;
      20'h08d2d: out <= 12'h666;
      20'h08d2e: out <= 12'hfff;
      20'h08d2f: out <= 12'h666;
      20'h08d30: out <= 12'hfff;
      20'h08d31: out <= 12'h666;
      20'h08d32: out <= 12'hfff;
      20'h08d33: out <= 12'h666;
      20'h08d34: out <= 12'hfff;
      20'h08d35: out <= 12'h666;
      20'h08d36: out <= 12'hfff;
      20'h08d37: out <= 12'h000;
      20'h08d38: out <= 12'h222;
      20'h08d39: out <= 12'h666;
      20'h08d3a: out <= 12'h666;
      20'h08d3b: out <= 12'hbbb;
      20'h08d3c: out <= 12'h666;
      20'h08d3d: out <= 12'h222;
      20'h08d3e: out <= 12'h222;
      20'h08d3f: out <= 12'hbbb;
      20'h08d40: out <= 12'hfff;
      20'h08d41: out <= 12'hbbb;
      20'h08d42: out <= 12'h222;
      20'h08d43: out <= 12'h222;
      20'h08d44: out <= 12'h666;
      20'h08d45: out <= 12'hbbb;
      20'h08d46: out <= 12'h666;
      20'h08d47: out <= 12'h666;
      20'h08d48: out <= 12'h000;
      20'h08d49: out <= 12'h666;
      20'h08d4a: out <= 12'hfff;
      20'h08d4b: out <= 12'hbbb;
      20'h08d4c: out <= 12'h666;
      20'h08d4d: out <= 12'h000;
      20'h08d4e: out <= 12'h000;
      20'h08d4f: out <= 12'hbbb;
      20'h08d50: out <= 12'hfff;
      20'h08d51: out <= 12'hbbb;
      20'h08d52: out <= 12'h000;
      20'h08d53: out <= 12'h000;
      20'h08d54: out <= 12'h666;
      20'h08d55: out <= 12'hbbb;
      20'h08d56: out <= 12'hfff;
      20'h08d57: out <= 12'h666;
      20'h08d58: out <= 12'h222;
      20'h08d59: out <= 12'h666;
      20'h08d5a: out <= 12'hfff;
      20'h08d5b: out <= 12'h666;
      20'h08d5c: out <= 12'hfff;
      20'h08d5d: out <= 12'h666;
      20'h08d5e: out <= 12'hfff;
      20'h08d5f: out <= 12'h666;
      20'h08d60: out <= 12'hfff;
      20'h08d61: out <= 12'h666;
      20'h08d62: out <= 12'hfff;
      20'h08d63: out <= 12'h666;
      20'h08d64: out <= 12'hfff;
      20'h08d65: out <= 12'h666;
      20'h08d66: out <= 12'hfff;
      20'h08d67: out <= 12'h222;
      20'h08d68: out <= 12'h000;
      20'h08d69: out <= 12'hfff;
      20'h08d6a: out <= 12'h666;
      20'h08d6b: out <= 12'hfff;
      20'h08d6c: out <= 12'h666;
      20'h08d6d: out <= 12'hfff;
      20'h08d6e: out <= 12'h666;
      20'h08d6f: out <= 12'hfff;
      20'h08d70: out <= 12'h666;
      20'h08d71: out <= 12'hfff;
      20'h08d72: out <= 12'h666;
      20'h08d73: out <= 12'hfff;
      20'h08d74: out <= 12'h666;
      20'h08d75: out <= 12'hfff;
      20'h08d76: out <= 12'h666;
      20'h08d77: out <= 12'h000;
      20'h08d78: out <= 12'h222;
      20'h08d79: out <= 12'h666;
      20'h08d7a: out <= 12'hfff;
      20'h08d7b: out <= 12'hbbb;
      20'h08d7c: out <= 12'h666;
      20'h08d7d: out <= 12'h222;
      20'h08d7e: out <= 12'h666;
      20'h08d7f: out <= 12'h666;
      20'h08d80: out <= 12'h666;
      20'h08d81: out <= 12'h666;
      20'h08d82: out <= 12'h666;
      20'h08d83: out <= 12'h222;
      20'h08d84: out <= 12'h666;
      20'h08d85: out <= 12'hbbb;
      20'h08d86: out <= 12'hfff;
      20'h08d87: out <= 12'h666;
      20'h08d88: out <= 12'h000;
      20'h08d89: out <= 12'h666;
      20'h08d8a: out <= 12'h666;
      20'h08d8b: out <= 12'hbbb;
      20'h08d8c: out <= 12'h666;
      20'h08d8d: out <= 12'h000;
      20'h08d8e: out <= 12'h666;
      20'h08d8f: out <= 12'h666;
      20'h08d90: out <= 12'h666;
      20'h08d91: out <= 12'h666;
      20'h08d92: out <= 12'h666;
      20'h08d93: out <= 12'h000;
      20'h08d94: out <= 12'h666;
      20'h08d95: out <= 12'hbbb;
      20'h08d96: out <= 12'h666;
      20'h08d97: out <= 12'h666;
      20'h08d98: out <= 12'h603;
      20'h08d99: out <= 12'h603;
      20'h08d9a: out <= 12'h603;
      20'h08d9b: out <= 12'h603;
      20'h08d9c: out <= 12'h603;
      20'h08d9d: out <= 12'h603;
      20'h08d9e: out <= 12'h603;
      20'h08d9f: out <= 12'h603;
      20'h08da0: out <= 12'h603;
      20'h08da1: out <= 12'h603;
      20'h08da2: out <= 12'h603;
      20'h08da3: out <= 12'h603;
      20'h08da4: out <= 12'h603;
      20'h08da5: out <= 12'h603;
      20'h08da6: out <= 12'h603;
      20'h08da7: out <= 12'h603;
      20'h08da8: out <= 12'h603;
      20'h08da9: out <= 12'h603;
      20'h08daa: out <= 12'h603;
      20'h08dab: out <= 12'h603;
      20'h08dac: out <= 12'h603;
      20'h08dad: out <= 12'h603;
      20'h08dae: out <= 12'h603;
      20'h08daf: out <= 12'h603;
      20'h08db0: out <= 12'h603;
      20'h08db1: out <= 12'h603;
      20'h08db2: out <= 12'h603;
      20'h08db3: out <= 12'h603;
      20'h08db4: out <= 12'h603;
      20'h08db5: out <= 12'h603;
      20'h08db6: out <= 12'h603;
      20'h08db7: out <= 12'h603;
      20'h08db8: out <= 12'h603;
      20'h08db9: out <= 12'h603;
      20'h08dba: out <= 12'h603;
      20'h08dbb: out <= 12'h603;
      20'h08dbc: out <= 12'h603;
      20'h08dbd: out <= 12'h603;
      20'h08dbe: out <= 12'h603;
      20'h08dbf: out <= 12'h603;
      20'h08dc0: out <= 12'h603;
      20'h08dc1: out <= 12'h603;
      20'h08dc2: out <= 12'h603;
      20'h08dc3: out <= 12'h603;
      20'h08dc4: out <= 12'h603;
      20'h08dc5: out <= 12'h603;
      20'h08dc6: out <= 12'h603;
      20'h08dc7: out <= 12'h603;
      20'h08dc8: out <= 12'h603;
      20'h08dc9: out <= 12'h603;
      20'h08dca: out <= 12'h603;
      20'h08dcb: out <= 12'h603;
      20'h08dcc: out <= 12'h603;
      20'h08dcd: out <= 12'h603;
      20'h08dce: out <= 12'h603;
      20'h08dcf: out <= 12'h603;
      20'h08dd0: out <= 12'h603;
      20'h08dd1: out <= 12'h603;
      20'h08dd2: out <= 12'h603;
      20'h08dd3: out <= 12'h603;
      20'h08dd4: out <= 12'h603;
      20'h08dd5: out <= 12'h603;
      20'h08dd6: out <= 12'h603;
      20'h08dd7: out <= 12'h603;
      20'h08dd8: out <= 12'h603;
      20'h08dd9: out <= 12'h603;
      20'h08dda: out <= 12'h603;
      20'h08ddb: out <= 12'h603;
      20'h08ddc: out <= 12'h603;
      20'h08ddd: out <= 12'h603;
      20'h08dde: out <= 12'h603;
      20'h08ddf: out <= 12'h603;
      20'h08de0: out <= 12'h603;
      20'h08de1: out <= 12'h603;
      20'h08de2: out <= 12'h603;
      20'h08de3: out <= 12'h603;
      20'h08de4: out <= 12'h603;
      20'h08de5: out <= 12'h603;
      20'h08de6: out <= 12'h603;
      20'h08de7: out <= 12'h603;
      20'h08de8: out <= 12'h603;
      20'h08de9: out <= 12'h603;
      20'h08dea: out <= 12'h603;
      20'h08deb: out <= 12'h603;
      20'h08dec: out <= 12'h603;
      20'h08ded: out <= 12'h603;
      20'h08dee: out <= 12'h603;
      20'h08def: out <= 12'h603;
      20'h08df0: out <= 12'hee9;
      20'h08df1: out <= 12'hf87;
      20'h08df2: out <= 12'hf87;
      20'h08df3: out <= 12'hf87;
      20'h08df4: out <= 12'hf87;
      20'h08df5: out <= 12'hf87;
      20'h08df6: out <= 12'hf87;
      20'h08df7: out <= 12'hb27;
      20'h08df8: out <= 12'h000;
      20'h08df9: out <= 12'h000;
      20'h08dfa: out <= 12'h000;
      20'h08dfb: out <= 12'h000;
      20'h08dfc: out <= 12'h000;
      20'h08dfd: out <= 12'h000;
      20'h08dfe: out <= 12'h000;
      20'h08dff: out <= 12'h000;
      20'h08e00: out <= 12'h8d0;
      20'h08e01: out <= 12'h8d0;
      20'h08e02: out <= 12'h000;
      20'h08e03: out <= 12'h000;
      20'h08e04: out <= 12'h000;
      20'h08e05: out <= 12'h8d0;
      20'h08e06: out <= 12'h8d0;
      20'h08e07: out <= 12'h000;
      20'h08e08: out <= 12'h8d0;
      20'h08e09: out <= 12'h8d0;
      20'h08e0a: out <= 12'h000;
      20'h08e0b: out <= 12'h000;
      20'h08e0c: out <= 12'h8d0;
      20'h08e0d: out <= 12'h8d0;
      20'h08e0e: out <= 12'h000;
      20'h08e0f: out <= 12'h8d0;
      20'h08e10: out <= 12'h8d0;
      20'h08e11: out <= 12'h000;
      20'h08e12: out <= 12'h000;
      20'h08e13: out <= 12'h000;
      20'h08e14: out <= 12'h000;
      20'h08e15: out <= 12'h8d0;
      20'h08e16: out <= 12'h8d0;
      20'h08e17: out <= 12'h8d0;
      20'h08e18: out <= 12'h8d0;
      20'h08e19: out <= 12'h8d0;
      20'h08e1a: out <= 12'h8d0;
      20'h08e1b: out <= 12'h000;
      20'h08e1c: out <= 12'h8d0;
      20'h08e1d: out <= 12'h8d0;
      20'h08e1e: out <= 12'h000;
      20'h08e1f: out <= 12'h000;
      20'h08e20: out <= 12'h000;
      20'h08e21: out <= 12'h8d0;
      20'h08e22: out <= 12'h8d0;
      20'h08e23: out <= 12'h000;
      20'h08e24: out <= 12'h000;
      20'h08e25: out <= 12'h000;
      20'h08e26: out <= 12'h000;
      20'h08e27: out <= 12'h000;
      20'h08e28: out <= 12'h000;
      20'h08e29: out <= 12'h000;
      20'h08e2a: out <= 12'h000;
      20'h08e2b: out <= 12'h000;
      20'h08e2c: out <= 12'h000;
      20'h08e2d: out <= 12'h000;
      20'h08e2e: out <= 12'h000;
      20'h08e2f: out <= 12'h000;
      20'h08e30: out <= 12'h222;
      20'h08e31: out <= 12'hbbb;
      20'h08e32: out <= 12'hbbb;
      20'h08e33: out <= 12'h666;
      20'h08e34: out <= 12'h666;
      20'h08e35: out <= 12'h666;
      20'h08e36: out <= 12'h666;
      20'h08e37: out <= 12'h666;
      20'h08e38: out <= 12'h666;
      20'h08e39: out <= 12'h666;
      20'h08e3a: out <= 12'h666;
      20'h08e3b: out <= 12'h666;
      20'h08e3c: out <= 12'hbbb;
      20'h08e3d: out <= 12'hbbb;
      20'h08e3e: out <= 12'hbbb;
      20'h08e3f: out <= 12'h222;
      20'h08e40: out <= 12'h000;
      20'h08e41: out <= 12'hbbb;
      20'h08e42: out <= 12'hbbb;
      20'h08e43: out <= 12'h666;
      20'h08e44: out <= 12'h666;
      20'h08e45: out <= 12'h666;
      20'h08e46: out <= 12'h666;
      20'h08e47: out <= 12'h666;
      20'h08e48: out <= 12'h666;
      20'h08e49: out <= 12'h666;
      20'h08e4a: out <= 12'h666;
      20'h08e4b: out <= 12'h666;
      20'h08e4c: out <= 12'hbbb;
      20'h08e4d: out <= 12'hbbb;
      20'h08e4e: out <= 12'hbbb;
      20'h08e4f: out <= 12'h000;
      20'h08e50: out <= 12'h222;
      20'h08e51: out <= 12'h666;
      20'h08e52: out <= 12'hfff;
      20'h08e53: out <= 12'hbbb;
      20'h08e54: out <= 12'h666;
      20'h08e55: out <= 12'h222;
      20'h08e56: out <= 12'h222;
      20'h08e57: out <= 12'hbbb;
      20'h08e58: out <= 12'hfff;
      20'h08e59: out <= 12'hbbb;
      20'h08e5a: out <= 12'h222;
      20'h08e5b: out <= 12'h222;
      20'h08e5c: out <= 12'h666;
      20'h08e5d: out <= 12'hbbb;
      20'h08e5e: out <= 12'hfff;
      20'h08e5f: out <= 12'h666;
      20'h08e60: out <= 12'h000;
      20'h08e61: out <= 12'h666;
      20'h08e62: out <= 12'h666;
      20'h08e63: out <= 12'hbbb;
      20'h08e64: out <= 12'h666;
      20'h08e65: out <= 12'h000;
      20'h08e66: out <= 12'h000;
      20'h08e67: out <= 12'hbbb;
      20'h08e68: out <= 12'hfff;
      20'h08e69: out <= 12'hbbb;
      20'h08e6a: out <= 12'h000;
      20'h08e6b: out <= 12'h000;
      20'h08e6c: out <= 12'h666;
      20'h08e6d: out <= 12'hbbb;
      20'h08e6e: out <= 12'h666;
      20'h08e6f: out <= 12'h666;
      20'h08e70: out <= 12'h222;
      20'h08e71: out <= 12'hbbb;
      20'h08e72: out <= 12'hbbb;
      20'h08e73: out <= 12'hbbb;
      20'h08e74: out <= 12'h666;
      20'h08e75: out <= 12'h666;
      20'h08e76: out <= 12'h666;
      20'h08e77: out <= 12'h666;
      20'h08e78: out <= 12'h666;
      20'h08e79: out <= 12'h666;
      20'h08e7a: out <= 12'h666;
      20'h08e7b: out <= 12'h666;
      20'h08e7c: out <= 12'h666;
      20'h08e7d: out <= 12'hbbb;
      20'h08e7e: out <= 12'hbbb;
      20'h08e7f: out <= 12'h222;
      20'h08e80: out <= 12'h000;
      20'h08e81: out <= 12'hbbb;
      20'h08e82: out <= 12'hbbb;
      20'h08e83: out <= 12'hbbb;
      20'h08e84: out <= 12'h666;
      20'h08e85: out <= 12'h666;
      20'h08e86: out <= 12'h666;
      20'h08e87: out <= 12'h666;
      20'h08e88: out <= 12'h666;
      20'h08e89: out <= 12'h666;
      20'h08e8a: out <= 12'h666;
      20'h08e8b: out <= 12'h666;
      20'h08e8c: out <= 12'h666;
      20'h08e8d: out <= 12'hbbb;
      20'h08e8e: out <= 12'hbbb;
      20'h08e8f: out <= 12'h000;
      20'h08e90: out <= 12'h222;
      20'h08e91: out <= 12'h666;
      20'h08e92: out <= 12'h666;
      20'h08e93: out <= 12'hbbb;
      20'h08e94: out <= 12'h666;
      20'h08e95: out <= 12'h666;
      20'h08e96: out <= 12'hfff;
      20'h08e97: out <= 12'hbbb;
      20'h08e98: out <= 12'h666;
      20'h08e99: out <= 12'hbbb;
      20'h08e9a: out <= 12'hfff;
      20'h08e9b: out <= 12'h666;
      20'h08e9c: out <= 12'h666;
      20'h08e9d: out <= 12'hbbb;
      20'h08e9e: out <= 12'h666;
      20'h08e9f: out <= 12'h666;
      20'h08ea0: out <= 12'h000;
      20'h08ea1: out <= 12'h666;
      20'h08ea2: out <= 12'hfff;
      20'h08ea3: out <= 12'hbbb;
      20'h08ea4: out <= 12'h666;
      20'h08ea5: out <= 12'h666;
      20'h08ea6: out <= 12'hfff;
      20'h08ea7: out <= 12'hbbb;
      20'h08ea8: out <= 12'h666;
      20'h08ea9: out <= 12'hbbb;
      20'h08eaa: out <= 12'hfff;
      20'h08eab: out <= 12'h666;
      20'h08eac: out <= 12'h666;
      20'h08ead: out <= 12'hbbb;
      20'h08eae: out <= 12'hfff;
      20'h08eaf: out <= 12'h666;
      20'h08eb0: out <= 12'h603;
      20'h08eb1: out <= 12'h603;
      20'h08eb2: out <= 12'h603;
      20'h08eb3: out <= 12'h603;
      20'h08eb4: out <= 12'h603;
      20'h08eb5: out <= 12'h603;
      20'h08eb6: out <= 12'h603;
      20'h08eb7: out <= 12'h603;
      20'h08eb8: out <= 12'h603;
      20'h08eb9: out <= 12'h603;
      20'h08eba: out <= 12'h603;
      20'h08ebb: out <= 12'h603;
      20'h08ebc: out <= 12'h603;
      20'h08ebd: out <= 12'h603;
      20'h08ebe: out <= 12'h603;
      20'h08ebf: out <= 12'h603;
      20'h08ec0: out <= 12'h603;
      20'h08ec1: out <= 12'h603;
      20'h08ec2: out <= 12'h603;
      20'h08ec3: out <= 12'h603;
      20'h08ec4: out <= 12'h603;
      20'h08ec5: out <= 12'h603;
      20'h08ec6: out <= 12'h603;
      20'h08ec7: out <= 12'h603;
      20'h08ec8: out <= 12'h603;
      20'h08ec9: out <= 12'h603;
      20'h08eca: out <= 12'h603;
      20'h08ecb: out <= 12'h603;
      20'h08ecc: out <= 12'h603;
      20'h08ecd: out <= 12'h603;
      20'h08ece: out <= 12'h603;
      20'h08ecf: out <= 12'h603;
      20'h08ed0: out <= 12'h603;
      20'h08ed1: out <= 12'h603;
      20'h08ed2: out <= 12'h603;
      20'h08ed3: out <= 12'h603;
      20'h08ed4: out <= 12'h603;
      20'h08ed5: out <= 12'h603;
      20'h08ed6: out <= 12'h603;
      20'h08ed7: out <= 12'h603;
      20'h08ed8: out <= 12'h603;
      20'h08ed9: out <= 12'h603;
      20'h08eda: out <= 12'h603;
      20'h08edb: out <= 12'h603;
      20'h08edc: out <= 12'h603;
      20'h08edd: out <= 12'h603;
      20'h08ede: out <= 12'h603;
      20'h08edf: out <= 12'h603;
      20'h08ee0: out <= 12'h603;
      20'h08ee1: out <= 12'h603;
      20'h08ee2: out <= 12'h603;
      20'h08ee3: out <= 12'h603;
      20'h08ee4: out <= 12'h603;
      20'h08ee5: out <= 12'h603;
      20'h08ee6: out <= 12'h603;
      20'h08ee7: out <= 12'h603;
      20'h08ee8: out <= 12'h603;
      20'h08ee9: out <= 12'h603;
      20'h08eea: out <= 12'h603;
      20'h08eeb: out <= 12'h603;
      20'h08eec: out <= 12'h603;
      20'h08eed: out <= 12'h603;
      20'h08eee: out <= 12'h603;
      20'h08eef: out <= 12'h603;
      20'h08ef0: out <= 12'h603;
      20'h08ef1: out <= 12'h603;
      20'h08ef2: out <= 12'h603;
      20'h08ef3: out <= 12'h603;
      20'h08ef4: out <= 12'h603;
      20'h08ef5: out <= 12'h603;
      20'h08ef6: out <= 12'h603;
      20'h08ef7: out <= 12'h603;
      20'h08ef8: out <= 12'h603;
      20'h08ef9: out <= 12'h603;
      20'h08efa: out <= 12'h603;
      20'h08efb: out <= 12'h603;
      20'h08efc: out <= 12'h603;
      20'h08efd: out <= 12'h603;
      20'h08efe: out <= 12'h603;
      20'h08eff: out <= 12'h603;
      20'h08f00: out <= 12'h603;
      20'h08f01: out <= 12'h603;
      20'h08f02: out <= 12'h603;
      20'h08f03: out <= 12'h603;
      20'h08f04: out <= 12'h603;
      20'h08f05: out <= 12'h603;
      20'h08f06: out <= 12'h603;
      20'h08f07: out <= 12'h603;
      20'h08f08: out <= 12'hee9;
      20'h08f09: out <= 12'hf87;
      20'h08f0a: out <= 12'hee9;
      20'h08f0b: out <= 12'hee9;
      20'h08f0c: out <= 12'hee9;
      20'h08f0d: out <= 12'hb27;
      20'h08f0e: out <= 12'hf87;
      20'h08f0f: out <= 12'hb27;
      20'h08f10: out <= 12'h000;
      20'h08f11: out <= 12'h000;
      20'h08f12: out <= 12'h000;
      20'h08f13: out <= 12'h000;
      20'h08f14: out <= 12'h000;
      20'h08f15: out <= 12'h000;
      20'h08f16: out <= 12'h000;
      20'h08f17: out <= 12'h000;
      20'h08f18: out <= 12'h000;
      20'h08f19: out <= 12'h000;
      20'h08f1a: out <= 12'h000;
      20'h08f1b: out <= 12'h000;
      20'h08f1c: out <= 12'h000;
      20'h08f1d: out <= 12'h8d0;
      20'h08f1e: out <= 12'h8d0;
      20'h08f1f: out <= 12'h000;
      20'h08f20: out <= 12'h8d0;
      20'h08f21: out <= 12'h8d0;
      20'h08f22: out <= 12'h000;
      20'h08f23: out <= 12'h000;
      20'h08f24: out <= 12'h8d0;
      20'h08f25: out <= 12'h8d0;
      20'h08f26: out <= 12'h000;
      20'h08f27: out <= 12'h8d0;
      20'h08f28: out <= 12'h8d0;
      20'h08f29: out <= 12'h000;
      20'h08f2a: out <= 12'h000;
      20'h08f2b: out <= 12'h000;
      20'h08f2c: out <= 12'h000;
      20'h08f2d: out <= 12'h8d0;
      20'h08f2e: out <= 12'h8d0;
      20'h08f2f: out <= 12'h000;
      20'h08f30: out <= 12'h000;
      20'h08f31: out <= 12'h8d0;
      20'h08f32: out <= 12'h8d0;
      20'h08f33: out <= 12'h000;
      20'h08f34: out <= 12'h8d0;
      20'h08f35: out <= 12'h8d0;
      20'h08f36: out <= 12'h000;
      20'h08f37: out <= 12'h000;
      20'h08f38: out <= 12'h000;
      20'h08f39: out <= 12'h8d0;
      20'h08f3a: out <= 12'h8d0;
      20'h08f3b: out <= 12'h000;
      20'h08f3c: out <= 12'h000;
      20'h08f3d: out <= 12'h000;
      20'h08f3e: out <= 12'h000;
      20'h08f3f: out <= 12'h000;
      20'h08f40: out <= 12'h000;
      20'h08f41: out <= 12'h000;
      20'h08f42: out <= 12'h000;
      20'h08f43: out <= 12'h000;
      20'h08f44: out <= 12'h000;
      20'h08f45: out <= 12'h000;
      20'h08f46: out <= 12'h000;
      20'h08f47: out <= 12'h000;
      20'h08f48: out <= 12'h222;
      20'h08f49: out <= 12'h666;
      20'h08f4a: out <= 12'h666;
      20'h08f4b: out <= 12'h666;
      20'h08f4c: out <= 12'hbbb;
      20'h08f4d: out <= 12'hbbb;
      20'h08f4e: out <= 12'hbbb;
      20'h08f4f: out <= 12'hbbb;
      20'h08f50: out <= 12'hbbb;
      20'h08f51: out <= 12'hbbb;
      20'h08f52: out <= 12'hbbb;
      20'h08f53: out <= 12'h666;
      20'h08f54: out <= 12'h666;
      20'h08f55: out <= 12'h666;
      20'h08f56: out <= 12'h666;
      20'h08f57: out <= 12'h222;
      20'h08f58: out <= 12'h000;
      20'h08f59: out <= 12'h666;
      20'h08f5a: out <= 12'h666;
      20'h08f5b: out <= 12'h666;
      20'h08f5c: out <= 12'hbbb;
      20'h08f5d: out <= 12'hbbb;
      20'h08f5e: out <= 12'hbbb;
      20'h08f5f: out <= 12'hbbb;
      20'h08f60: out <= 12'hbbb;
      20'h08f61: out <= 12'hbbb;
      20'h08f62: out <= 12'hbbb;
      20'h08f63: out <= 12'h666;
      20'h08f64: out <= 12'h666;
      20'h08f65: out <= 12'h666;
      20'h08f66: out <= 12'h666;
      20'h08f67: out <= 12'h000;
      20'h08f68: out <= 12'h222;
      20'h08f69: out <= 12'h666;
      20'h08f6a: out <= 12'h666;
      20'h08f6b: out <= 12'hbbb;
      20'h08f6c: out <= 12'h666;
      20'h08f6d: out <= 12'h666;
      20'h08f6e: out <= 12'h666;
      20'h08f6f: out <= 12'hbbb;
      20'h08f70: out <= 12'hfff;
      20'h08f71: out <= 12'hbbb;
      20'h08f72: out <= 12'h666;
      20'h08f73: out <= 12'h666;
      20'h08f74: out <= 12'h666;
      20'h08f75: out <= 12'hbbb;
      20'h08f76: out <= 12'h666;
      20'h08f77: out <= 12'h666;
      20'h08f78: out <= 12'h000;
      20'h08f79: out <= 12'h666;
      20'h08f7a: out <= 12'hfff;
      20'h08f7b: out <= 12'hbbb;
      20'h08f7c: out <= 12'h666;
      20'h08f7d: out <= 12'h666;
      20'h08f7e: out <= 12'h666;
      20'h08f7f: out <= 12'hbbb;
      20'h08f80: out <= 12'hfff;
      20'h08f81: out <= 12'hbbb;
      20'h08f82: out <= 12'h666;
      20'h08f83: out <= 12'h666;
      20'h08f84: out <= 12'h666;
      20'h08f85: out <= 12'hbbb;
      20'h08f86: out <= 12'hfff;
      20'h08f87: out <= 12'h666;
      20'h08f88: out <= 12'h222;
      20'h08f89: out <= 12'h666;
      20'h08f8a: out <= 12'h666;
      20'h08f8b: out <= 12'h666;
      20'h08f8c: out <= 12'h666;
      20'h08f8d: out <= 12'hbbb;
      20'h08f8e: out <= 12'hbbb;
      20'h08f8f: out <= 12'hbbb;
      20'h08f90: out <= 12'hbbb;
      20'h08f91: out <= 12'hbbb;
      20'h08f92: out <= 12'hbbb;
      20'h08f93: out <= 12'hbbb;
      20'h08f94: out <= 12'h666;
      20'h08f95: out <= 12'h666;
      20'h08f96: out <= 12'h666;
      20'h08f97: out <= 12'h222;
      20'h08f98: out <= 12'h000;
      20'h08f99: out <= 12'h666;
      20'h08f9a: out <= 12'h666;
      20'h08f9b: out <= 12'h666;
      20'h08f9c: out <= 12'h666;
      20'h08f9d: out <= 12'hbbb;
      20'h08f9e: out <= 12'hbbb;
      20'h08f9f: out <= 12'hbbb;
      20'h08fa0: out <= 12'hbbb;
      20'h08fa1: out <= 12'hbbb;
      20'h08fa2: out <= 12'hbbb;
      20'h08fa3: out <= 12'hbbb;
      20'h08fa4: out <= 12'h666;
      20'h08fa5: out <= 12'h666;
      20'h08fa6: out <= 12'h666;
      20'h08fa7: out <= 12'h000;
      20'h08fa8: out <= 12'h222;
      20'h08fa9: out <= 12'h666;
      20'h08faa: out <= 12'hfff;
      20'h08fab: out <= 12'h666;
      20'h08fac: out <= 12'h666;
      20'h08fad: out <= 12'hfff;
      20'h08fae: out <= 12'h666;
      20'h08faf: out <= 12'h666;
      20'h08fb0: out <= 12'h666;
      20'h08fb1: out <= 12'h666;
      20'h08fb2: out <= 12'h666;
      20'h08fb3: out <= 12'hfff;
      20'h08fb4: out <= 12'h666;
      20'h08fb5: out <= 12'h666;
      20'h08fb6: out <= 12'hfff;
      20'h08fb7: out <= 12'h666;
      20'h08fb8: out <= 12'h000;
      20'h08fb9: out <= 12'h666;
      20'h08fba: out <= 12'h666;
      20'h08fbb: out <= 12'h666;
      20'h08fbc: out <= 12'h666;
      20'h08fbd: out <= 12'hfff;
      20'h08fbe: out <= 12'h666;
      20'h08fbf: out <= 12'h666;
      20'h08fc0: out <= 12'h666;
      20'h08fc1: out <= 12'h666;
      20'h08fc2: out <= 12'h666;
      20'h08fc3: out <= 12'hfff;
      20'h08fc4: out <= 12'h666;
      20'h08fc5: out <= 12'h666;
      20'h08fc6: out <= 12'h666;
      20'h08fc7: out <= 12'h666;
      20'h08fc8: out <= 12'h603;
      20'h08fc9: out <= 12'h603;
      20'h08fca: out <= 12'h603;
      20'h08fcb: out <= 12'h603;
      20'h08fcc: out <= 12'h603;
      20'h08fcd: out <= 12'h603;
      20'h08fce: out <= 12'h603;
      20'h08fcf: out <= 12'h603;
      20'h08fd0: out <= 12'h603;
      20'h08fd1: out <= 12'h603;
      20'h08fd2: out <= 12'h603;
      20'h08fd3: out <= 12'h603;
      20'h08fd4: out <= 12'h603;
      20'h08fd5: out <= 12'h603;
      20'h08fd6: out <= 12'h603;
      20'h08fd7: out <= 12'h603;
      20'h08fd8: out <= 12'h603;
      20'h08fd9: out <= 12'h603;
      20'h08fda: out <= 12'h603;
      20'h08fdb: out <= 12'h603;
      20'h08fdc: out <= 12'h603;
      20'h08fdd: out <= 12'h603;
      20'h08fde: out <= 12'h603;
      20'h08fdf: out <= 12'h603;
      20'h08fe0: out <= 12'h603;
      20'h08fe1: out <= 12'h603;
      20'h08fe2: out <= 12'h603;
      20'h08fe3: out <= 12'h603;
      20'h08fe4: out <= 12'h603;
      20'h08fe5: out <= 12'h603;
      20'h08fe6: out <= 12'h603;
      20'h08fe7: out <= 12'h603;
      20'h08fe8: out <= 12'h603;
      20'h08fe9: out <= 12'h603;
      20'h08fea: out <= 12'h603;
      20'h08feb: out <= 12'h603;
      20'h08fec: out <= 12'h603;
      20'h08fed: out <= 12'h603;
      20'h08fee: out <= 12'h603;
      20'h08fef: out <= 12'h603;
      20'h08ff0: out <= 12'h603;
      20'h08ff1: out <= 12'h603;
      20'h08ff2: out <= 12'h603;
      20'h08ff3: out <= 12'h603;
      20'h08ff4: out <= 12'h603;
      20'h08ff5: out <= 12'h603;
      20'h08ff6: out <= 12'h603;
      20'h08ff7: out <= 12'h603;
      20'h08ff8: out <= 12'h603;
      20'h08ff9: out <= 12'h603;
      20'h08ffa: out <= 12'h603;
      20'h08ffb: out <= 12'h603;
      20'h08ffc: out <= 12'h603;
      20'h08ffd: out <= 12'h603;
      20'h08ffe: out <= 12'h603;
      20'h08fff: out <= 12'h603;
      20'h09000: out <= 12'h603;
      20'h09001: out <= 12'h603;
      20'h09002: out <= 12'h603;
      20'h09003: out <= 12'h603;
      20'h09004: out <= 12'h603;
      20'h09005: out <= 12'h603;
      20'h09006: out <= 12'h603;
      20'h09007: out <= 12'h603;
      20'h09008: out <= 12'h603;
      20'h09009: out <= 12'h603;
      20'h0900a: out <= 12'h603;
      20'h0900b: out <= 12'h603;
      20'h0900c: out <= 12'h603;
      20'h0900d: out <= 12'h603;
      20'h0900e: out <= 12'h603;
      20'h0900f: out <= 12'h603;
      20'h09010: out <= 12'h603;
      20'h09011: out <= 12'h603;
      20'h09012: out <= 12'h603;
      20'h09013: out <= 12'h603;
      20'h09014: out <= 12'h603;
      20'h09015: out <= 12'h603;
      20'h09016: out <= 12'h603;
      20'h09017: out <= 12'h603;
      20'h09018: out <= 12'h603;
      20'h09019: out <= 12'h603;
      20'h0901a: out <= 12'h603;
      20'h0901b: out <= 12'h603;
      20'h0901c: out <= 12'h603;
      20'h0901d: out <= 12'h603;
      20'h0901e: out <= 12'h603;
      20'h0901f: out <= 12'h603;
      20'h09020: out <= 12'hee9;
      20'h09021: out <= 12'hf87;
      20'h09022: out <= 12'hee9;
      20'h09023: out <= 12'hf87;
      20'h09024: out <= 12'hf87;
      20'h09025: out <= 12'hb27;
      20'h09026: out <= 12'hf87;
      20'h09027: out <= 12'hb27;
      20'h09028: out <= 12'h000;
      20'h09029: out <= 12'h000;
      20'h0902a: out <= 12'h000;
      20'h0902b: out <= 12'h000;
      20'h0902c: out <= 12'h000;
      20'h0902d: out <= 12'h000;
      20'h0902e: out <= 12'h000;
      20'h0902f: out <= 12'h000;
      20'h09030: out <= 12'h000;
      20'h09031: out <= 12'h000;
      20'h09032: out <= 12'h000;
      20'h09033: out <= 12'h8d0;
      20'h09034: out <= 12'h8d0;
      20'h09035: out <= 12'h8d0;
      20'h09036: out <= 12'h000;
      20'h09037: out <= 12'h000;
      20'h09038: out <= 12'h8d0;
      20'h09039: out <= 12'h8d0;
      20'h0903a: out <= 12'h8d0;
      20'h0903b: out <= 12'h8d0;
      20'h0903c: out <= 12'h8d0;
      20'h0903d: out <= 12'h000;
      20'h0903e: out <= 12'h000;
      20'h0903f: out <= 12'h8d0;
      20'h09040: out <= 12'h8d0;
      20'h09041: out <= 12'h000;
      20'h09042: out <= 12'h000;
      20'h09043: out <= 12'h000;
      20'h09044: out <= 12'h000;
      20'h09045: out <= 12'h8d0;
      20'h09046: out <= 12'h8d0;
      20'h09047: out <= 12'h000;
      20'h09048: out <= 12'h000;
      20'h09049: out <= 12'h8d0;
      20'h0904a: out <= 12'h8d0;
      20'h0904b: out <= 12'h000;
      20'h0904c: out <= 12'h000;
      20'h0904d: out <= 12'h8d0;
      20'h0904e: out <= 12'h8d0;
      20'h0904f: out <= 12'h8d0;
      20'h09050: out <= 12'h8d0;
      20'h09051: out <= 12'h8d0;
      20'h09052: out <= 12'h000;
      20'h09053: out <= 12'h000;
      20'h09054: out <= 12'h000;
      20'h09055: out <= 12'h000;
      20'h09056: out <= 12'h000;
      20'h09057: out <= 12'h000;
      20'h09058: out <= 12'h000;
      20'h09059: out <= 12'h000;
      20'h0905a: out <= 12'h000;
      20'h0905b: out <= 12'h000;
      20'h0905c: out <= 12'h000;
      20'h0905d: out <= 12'h000;
      20'h0905e: out <= 12'h000;
      20'h0905f: out <= 12'h000;
      20'h09060: out <= 12'h222;
      20'h09061: out <= 12'h222;
      20'h09062: out <= 12'h666;
      20'h09063: out <= 12'hfff;
      20'h09064: out <= 12'hfff;
      20'h09065: out <= 12'hbbb;
      20'h09066: out <= 12'h666;
      20'h09067: out <= 12'hbbb;
      20'h09068: out <= 12'h666;
      20'h09069: out <= 12'hbbb;
      20'h0906a: out <= 12'hfff;
      20'h0906b: out <= 12'hfff;
      20'h0906c: out <= 12'h666;
      20'h0906d: out <= 12'h222;
      20'h0906e: out <= 12'h222;
      20'h0906f: out <= 12'h222;
      20'h09070: out <= 12'h000;
      20'h09071: out <= 12'h000;
      20'h09072: out <= 12'h666;
      20'h09073: out <= 12'hfff;
      20'h09074: out <= 12'hfff;
      20'h09075: out <= 12'hbbb;
      20'h09076: out <= 12'h666;
      20'h09077: out <= 12'hbbb;
      20'h09078: out <= 12'h666;
      20'h09079: out <= 12'hbbb;
      20'h0907a: out <= 12'hfff;
      20'h0907b: out <= 12'hfff;
      20'h0907c: out <= 12'h666;
      20'h0907d: out <= 12'h000;
      20'h0907e: out <= 12'h000;
      20'h0907f: out <= 12'h000;
      20'h09080: out <= 12'h222;
      20'h09081: out <= 12'h666;
      20'h09082: out <= 12'hfff;
      20'h09083: out <= 12'h666;
      20'h09084: out <= 12'h666;
      20'h09085: out <= 12'hfff;
      20'h09086: out <= 12'h666;
      20'h09087: out <= 12'hbbb;
      20'h09088: out <= 12'hfff;
      20'h09089: out <= 12'hbbb;
      20'h0908a: out <= 12'h666;
      20'h0908b: out <= 12'hfff;
      20'h0908c: out <= 12'h666;
      20'h0908d: out <= 12'h666;
      20'h0908e: out <= 12'hfff;
      20'h0908f: out <= 12'h666;
      20'h09090: out <= 12'h000;
      20'h09091: out <= 12'h666;
      20'h09092: out <= 12'h666;
      20'h09093: out <= 12'h666;
      20'h09094: out <= 12'h666;
      20'h09095: out <= 12'hfff;
      20'h09096: out <= 12'h666;
      20'h09097: out <= 12'hbbb;
      20'h09098: out <= 12'hfff;
      20'h09099: out <= 12'hbbb;
      20'h0909a: out <= 12'h666;
      20'h0909b: out <= 12'hfff;
      20'h0909c: out <= 12'h666;
      20'h0909d: out <= 12'h666;
      20'h0909e: out <= 12'h666;
      20'h0909f: out <= 12'h666;
      20'h090a0: out <= 12'h222;
      20'h090a1: out <= 12'h222;
      20'h090a2: out <= 12'h222;
      20'h090a3: out <= 12'h666;
      20'h090a4: out <= 12'hfff;
      20'h090a5: out <= 12'hfff;
      20'h090a6: out <= 12'hbbb;
      20'h090a7: out <= 12'h666;
      20'h090a8: out <= 12'hbbb;
      20'h090a9: out <= 12'h666;
      20'h090aa: out <= 12'hbbb;
      20'h090ab: out <= 12'hfff;
      20'h090ac: out <= 12'hfff;
      20'h090ad: out <= 12'h666;
      20'h090ae: out <= 12'h222;
      20'h090af: out <= 12'h222;
      20'h090b0: out <= 12'h000;
      20'h090b1: out <= 12'h000;
      20'h090b2: out <= 12'h000;
      20'h090b3: out <= 12'h666;
      20'h090b4: out <= 12'hfff;
      20'h090b5: out <= 12'hfff;
      20'h090b6: out <= 12'hbbb;
      20'h090b7: out <= 12'h666;
      20'h090b8: out <= 12'hbbb;
      20'h090b9: out <= 12'h666;
      20'h090ba: out <= 12'hbbb;
      20'h090bb: out <= 12'hfff;
      20'h090bc: out <= 12'hfff;
      20'h090bd: out <= 12'h666;
      20'h090be: out <= 12'h000;
      20'h090bf: out <= 12'h000;
      20'h090c0: out <= 12'h222;
      20'h090c1: out <= 12'h666;
      20'h090c2: out <= 12'h666;
      20'h090c3: out <= 12'h666;
      20'h090c4: out <= 12'hbbb;
      20'h090c5: out <= 12'hfff;
      20'h090c6: out <= 12'h666;
      20'h090c7: out <= 12'hfff;
      20'h090c8: out <= 12'hfff;
      20'h090c9: out <= 12'hfff;
      20'h090ca: out <= 12'h666;
      20'h090cb: out <= 12'hfff;
      20'h090cc: out <= 12'hbbb;
      20'h090cd: out <= 12'h666;
      20'h090ce: out <= 12'h666;
      20'h090cf: out <= 12'h666;
      20'h090d0: out <= 12'h000;
      20'h090d1: out <= 12'h666;
      20'h090d2: out <= 12'hfff;
      20'h090d3: out <= 12'h666;
      20'h090d4: out <= 12'hbbb;
      20'h090d5: out <= 12'hfff;
      20'h090d6: out <= 12'h666;
      20'h090d7: out <= 12'hbbb;
      20'h090d8: out <= 12'hfff;
      20'h090d9: out <= 12'hfff;
      20'h090da: out <= 12'h666;
      20'h090db: out <= 12'hfff;
      20'h090dc: out <= 12'hbbb;
      20'h090dd: out <= 12'h666;
      20'h090de: out <= 12'hfff;
      20'h090df: out <= 12'h666;
      20'h090e0: out <= 12'h603;
      20'h090e1: out <= 12'h603;
      20'h090e2: out <= 12'h603;
      20'h090e3: out <= 12'h603;
      20'h090e4: out <= 12'h603;
      20'h090e5: out <= 12'h603;
      20'h090e6: out <= 12'h603;
      20'h090e7: out <= 12'h603;
      20'h090e8: out <= 12'h603;
      20'h090e9: out <= 12'h603;
      20'h090ea: out <= 12'h603;
      20'h090eb: out <= 12'h603;
      20'h090ec: out <= 12'h603;
      20'h090ed: out <= 12'h603;
      20'h090ee: out <= 12'h603;
      20'h090ef: out <= 12'h603;
      20'h090f0: out <= 12'h603;
      20'h090f1: out <= 12'h603;
      20'h090f2: out <= 12'h603;
      20'h090f3: out <= 12'h603;
      20'h090f4: out <= 12'h603;
      20'h090f5: out <= 12'h603;
      20'h090f6: out <= 12'h603;
      20'h090f7: out <= 12'h603;
      20'h090f8: out <= 12'h603;
      20'h090f9: out <= 12'h603;
      20'h090fa: out <= 12'h603;
      20'h090fb: out <= 12'h603;
      20'h090fc: out <= 12'h603;
      20'h090fd: out <= 12'h603;
      20'h090fe: out <= 12'h603;
      20'h090ff: out <= 12'h603;
      20'h09100: out <= 12'h603;
      20'h09101: out <= 12'h603;
      20'h09102: out <= 12'h603;
      20'h09103: out <= 12'h603;
      20'h09104: out <= 12'h603;
      20'h09105: out <= 12'h603;
      20'h09106: out <= 12'h603;
      20'h09107: out <= 12'h603;
      20'h09108: out <= 12'h603;
      20'h09109: out <= 12'h603;
      20'h0910a: out <= 12'h603;
      20'h0910b: out <= 12'h603;
      20'h0910c: out <= 12'h603;
      20'h0910d: out <= 12'h603;
      20'h0910e: out <= 12'h603;
      20'h0910f: out <= 12'h603;
      20'h09110: out <= 12'h603;
      20'h09111: out <= 12'h603;
      20'h09112: out <= 12'h603;
      20'h09113: out <= 12'h603;
      20'h09114: out <= 12'h603;
      20'h09115: out <= 12'h603;
      20'h09116: out <= 12'h603;
      20'h09117: out <= 12'h603;
      20'h09118: out <= 12'h603;
      20'h09119: out <= 12'h603;
      20'h0911a: out <= 12'h603;
      20'h0911b: out <= 12'h603;
      20'h0911c: out <= 12'h603;
      20'h0911d: out <= 12'h603;
      20'h0911e: out <= 12'h603;
      20'h0911f: out <= 12'h603;
      20'h09120: out <= 12'h603;
      20'h09121: out <= 12'h603;
      20'h09122: out <= 12'h603;
      20'h09123: out <= 12'h603;
      20'h09124: out <= 12'h603;
      20'h09125: out <= 12'h603;
      20'h09126: out <= 12'h603;
      20'h09127: out <= 12'h603;
      20'h09128: out <= 12'h603;
      20'h09129: out <= 12'h603;
      20'h0912a: out <= 12'h603;
      20'h0912b: out <= 12'h603;
      20'h0912c: out <= 12'h603;
      20'h0912d: out <= 12'h603;
      20'h0912e: out <= 12'h603;
      20'h0912f: out <= 12'h603;
      20'h09130: out <= 12'h603;
      20'h09131: out <= 12'h603;
      20'h09132: out <= 12'h603;
      20'h09133: out <= 12'h603;
      20'h09134: out <= 12'h603;
      20'h09135: out <= 12'h603;
      20'h09136: out <= 12'h603;
      20'h09137: out <= 12'h603;
      20'h09138: out <= 12'hee9;
      20'h09139: out <= 12'hf87;
      20'h0913a: out <= 12'hee9;
      20'h0913b: out <= 12'hf87;
      20'h0913c: out <= 12'hf87;
      20'h0913d: out <= 12'hb27;
      20'h0913e: out <= 12'hf87;
      20'h0913f: out <= 12'hb27;
      20'h09140: out <= 12'h000;
      20'h09141: out <= 12'h000;
      20'h09142: out <= 12'h000;
      20'h09143: out <= 12'h000;
      20'h09144: out <= 12'h000;
      20'h09145: out <= 12'h000;
      20'h09146: out <= 12'h000;
      20'h09147: out <= 12'h000;
      20'h09148: out <= 12'h000;
      20'h09149: out <= 12'h8d0;
      20'h0914a: out <= 12'h8d0;
      20'h0914b: out <= 12'h8d0;
      20'h0914c: out <= 12'h000;
      20'h0914d: out <= 12'h000;
      20'h0914e: out <= 12'h000;
      20'h0914f: out <= 12'h000;
      20'h09150: out <= 12'h8d0;
      20'h09151: out <= 12'h8d0;
      20'h09152: out <= 12'h000;
      20'h09153: out <= 12'h000;
      20'h09154: out <= 12'h000;
      20'h09155: out <= 12'h000;
      20'h09156: out <= 12'h000;
      20'h09157: out <= 12'h8d0;
      20'h09158: out <= 12'h8d0;
      20'h09159: out <= 12'h000;
      20'h0915a: out <= 12'h000;
      20'h0915b: out <= 12'h000;
      20'h0915c: out <= 12'h000;
      20'h0915d: out <= 12'h8d0;
      20'h0915e: out <= 12'h8d0;
      20'h0915f: out <= 12'h8d0;
      20'h09160: out <= 12'h8d0;
      20'h09161: out <= 12'h8d0;
      20'h09162: out <= 12'h8d0;
      20'h09163: out <= 12'h000;
      20'h09164: out <= 12'h000;
      20'h09165: out <= 12'h000;
      20'h09166: out <= 12'h8d0;
      20'h09167: out <= 12'h8d0;
      20'h09168: out <= 12'h8d0;
      20'h09169: out <= 12'h000;
      20'h0916a: out <= 12'h000;
      20'h0916b: out <= 12'h000;
      20'h0916c: out <= 12'h000;
      20'h0916d: out <= 12'h000;
      20'h0916e: out <= 12'h000;
      20'h0916f: out <= 12'h000;
      20'h09170: out <= 12'h000;
      20'h09171: out <= 12'h000;
      20'h09172: out <= 12'h000;
      20'h09173: out <= 12'h000;
      20'h09174: out <= 12'h000;
      20'h09175: out <= 12'h000;
      20'h09176: out <= 12'h000;
      20'h09177: out <= 12'h000;
      20'h09178: out <= 12'h222;
      20'h09179: out <= 12'h666;
      20'h0917a: out <= 12'hfff;
      20'h0917b: out <= 12'h666;
      20'h0917c: out <= 12'h666;
      20'h0917d: out <= 12'h666;
      20'h0917e: out <= 12'h666;
      20'h0917f: out <= 12'h666;
      20'h09180: out <= 12'h666;
      20'h09181: out <= 12'h666;
      20'h09182: out <= 12'h666;
      20'h09183: out <= 12'h666;
      20'h09184: out <= 12'h666;
      20'h09185: out <= 12'h222;
      20'h09186: out <= 12'h222;
      20'h09187: out <= 12'hbbb;
      20'h09188: out <= 12'h000;
      20'h09189: out <= 12'h666;
      20'h0918a: out <= 12'hfff;
      20'h0918b: out <= 12'h666;
      20'h0918c: out <= 12'h666;
      20'h0918d: out <= 12'h666;
      20'h0918e: out <= 12'h666;
      20'h0918f: out <= 12'h666;
      20'h09190: out <= 12'h666;
      20'h09191: out <= 12'h666;
      20'h09192: out <= 12'h666;
      20'h09193: out <= 12'h666;
      20'h09194: out <= 12'h666;
      20'h09195: out <= 12'h000;
      20'h09196: out <= 12'h000;
      20'h09197: out <= 12'hbbb;
      20'h09198: out <= 12'h222;
      20'h09199: out <= 12'h666;
      20'h0919a: out <= 12'h666;
      20'h0919b: out <= 12'h666;
      20'h0919c: out <= 12'hbbb;
      20'h0919d: out <= 12'hfff;
      20'h0919e: out <= 12'h666;
      20'h0919f: out <= 12'h666;
      20'h091a0: out <= 12'h666;
      20'h091a1: out <= 12'h666;
      20'h091a2: out <= 12'h666;
      20'h091a3: out <= 12'hfff;
      20'h091a4: out <= 12'hbbb;
      20'h091a5: out <= 12'h666;
      20'h091a6: out <= 12'h666;
      20'h091a7: out <= 12'h666;
      20'h091a8: out <= 12'h000;
      20'h091a9: out <= 12'h666;
      20'h091aa: out <= 12'hfff;
      20'h091ab: out <= 12'h666;
      20'h091ac: out <= 12'hbbb;
      20'h091ad: out <= 12'hfff;
      20'h091ae: out <= 12'h666;
      20'h091af: out <= 12'h666;
      20'h091b0: out <= 12'h666;
      20'h091b1: out <= 12'h666;
      20'h091b2: out <= 12'h666;
      20'h091b3: out <= 12'hfff;
      20'h091b4: out <= 12'hbbb;
      20'h091b5: out <= 12'h666;
      20'h091b6: out <= 12'hfff;
      20'h091b7: out <= 12'h666;
      20'h091b8: out <= 12'hbbb;
      20'h091b9: out <= 12'h222;
      20'h091ba: out <= 12'h222;
      20'h091bb: out <= 12'h666;
      20'h091bc: out <= 12'h666;
      20'h091bd: out <= 12'h666;
      20'h091be: out <= 12'h666;
      20'h091bf: out <= 12'h666;
      20'h091c0: out <= 12'h666;
      20'h091c1: out <= 12'h666;
      20'h091c2: out <= 12'h666;
      20'h091c3: out <= 12'h666;
      20'h091c4: out <= 12'h666;
      20'h091c5: out <= 12'hfff;
      20'h091c6: out <= 12'h666;
      20'h091c7: out <= 12'h222;
      20'h091c8: out <= 12'hbbb;
      20'h091c9: out <= 12'h000;
      20'h091ca: out <= 12'h000;
      20'h091cb: out <= 12'h666;
      20'h091cc: out <= 12'h666;
      20'h091cd: out <= 12'h666;
      20'h091ce: out <= 12'h666;
      20'h091cf: out <= 12'h666;
      20'h091d0: out <= 12'h666;
      20'h091d1: out <= 12'h666;
      20'h091d2: out <= 12'h666;
      20'h091d3: out <= 12'h666;
      20'h091d4: out <= 12'h666;
      20'h091d5: out <= 12'hfff;
      20'h091d6: out <= 12'h666;
      20'h091d7: out <= 12'h000;
      20'h091d8: out <= 12'h222;
      20'h091d9: out <= 12'h666;
      20'h091da: out <= 12'hfff;
      20'h091db: out <= 12'h666;
      20'h091dc: out <= 12'hbbb;
      20'h091dd: out <= 12'hbbb;
      20'h091de: out <= 12'h666;
      20'h091df: out <= 12'hbbb;
      20'h091e0: out <= 12'hfff;
      20'h091e1: out <= 12'hfff;
      20'h091e2: out <= 12'h666;
      20'h091e3: out <= 12'hbbb;
      20'h091e4: out <= 12'hbbb;
      20'h091e5: out <= 12'h666;
      20'h091e6: out <= 12'hfff;
      20'h091e7: out <= 12'h666;
      20'h091e8: out <= 12'h000;
      20'h091e9: out <= 12'h666;
      20'h091ea: out <= 12'h666;
      20'h091eb: out <= 12'h666;
      20'h091ec: out <= 12'hbbb;
      20'h091ed: out <= 12'hbbb;
      20'h091ee: out <= 12'h666;
      20'h091ef: out <= 12'hbbb;
      20'h091f0: out <= 12'hbbb;
      20'h091f1: out <= 12'hfff;
      20'h091f2: out <= 12'h666;
      20'h091f3: out <= 12'hbbb;
      20'h091f4: out <= 12'hbbb;
      20'h091f5: out <= 12'h666;
      20'h091f6: out <= 12'h666;
      20'h091f7: out <= 12'h666;
      20'h091f8: out <= 12'h603;
      20'h091f9: out <= 12'h603;
      20'h091fa: out <= 12'h603;
      20'h091fb: out <= 12'h603;
      20'h091fc: out <= 12'h603;
      20'h091fd: out <= 12'h603;
      20'h091fe: out <= 12'h603;
      20'h091ff: out <= 12'h603;
      20'h09200: out <= 12'h603;
      20'h09201: out <= 12'h603;
      20'h09202: out <= 12'h603;
      20'h09203: out <= 12'h603;
      20'h09204: out <= 12'h603;
      20'h09205: out <= 12'h603;
      20'h09206: out <= 12'h603;
      20'h09207: out <= 12'h603;
      20'h09208: out <= 12'h603;
      20'h09209: out <= 12'h603;
      20'h0920a: out <= 12'h603;
      20'h0920b: out <= 12'h603;
      20'h0920c: out <= 12'h603;
      20'h0920d: out <= 12'h603;
      20'h0920e: out <= 12'h603;
      20'h0920f: out <= 12'h603;
      20'h09210: out <= 12'h603;
      20'h09211: out <= 12'h603;
      20'h09212: out <= 12'h603;
      20'h09213: out <= 12'h603;
      20'h09214: out <= 12'h603;
      20'h09215: out <= 12'h603;
      20'h09216: out <= 12'h603;
      20'h09217: out <= 12'h603;
      20'h09218: out <= 12'h603;
      20'h09219: out <= 12'h603;
      20'h0921a: out <= 12'h603;
      20'h0921b: out <= 12'h603;
      20'h0921c: out <= 12'h603;
      20'h0921d: out <= 12'h603;
      20'h0921e: out <= 12'h603;
      20'h0921f: out <= 12'h603;
      20'h09220: out <= 12'h603;
      20'h09221: out <= 12'h603;
      20'h09222: out <= 12'h603;
      20'h09223: out <= 12'h603;
      20'h09224: out <= 12'h603;
      20'h09225: out <= 12'h603;
      20'h09226: out <= 12'h603;
      20'h09227: out <= 12'h603;
      20'h09228: out <= 12'h603;
      20'h09229: out <= 12'h603;
      20'h0922a: out <= 12'h603;
      20'h0922b: out <= 12'h603;
      20'h0922c: out <= 12'h603;
      20'h0922d: out <= 12'h603;
      20'h0922e: out <= 12'h603;
      20'h0922f: out <= 12'h603;
      20'h09230: out <= 12'h603;
      20'h09231: out <= 12'h603;
      20'h09232: out <= 12'h603;
      20'h09233: out <= 12'h603;
      20'h09234: out <= 12'h603;
      20'h09235: out <= 12'h603;
      20'h09236: out <= 12'h603;
      20'h09237: out <= 12'h603;
      20'h09238: out <= 12'h603;
      20'h09239: out <= 12'h603;
      20'h0923a: out <= 12'h603;
      20'h0923b: out <= 12'h603;
      20'h0923c: out <= 12'h603;
      20'h0923d: out <= 12'h603;
      20'h0923e: out <= 12'h603;
      20'h0923f: out <= 12'h603;
      20'h09240: out <= 12'h603;
      20'h09241: out <= 12'h603;
      20'h09242: out <= 12'h603;
      20'h09243: out <= 12'h603;
      20'h09244: out <= 12'h603;
      20'h09245: out <= 12'h603;
      20'h09246: out <= 12'h603;
      20'h09247: out <= 12'h603;
      20'h09248: out <= 12'h603;
      20'h09249: out <= 12'h603;
      20'h0924a: out <= 12'h603;
      20'h0924b: out <= 12'h603;
      20'h0924c: out <= 12'h603;
      20'h0924d: out <= 12'h603;
      20'h0924e: out <= 12'h603;
      20'h0924f: out <= 12'h603;
      20'h09250: out <= 12'hee9;
      20'h09251: out <= 12'hf87;
      20'h09252: out <= 12'hee9;
      20'h09253: out <= 12'hb27;
      20'h09254: out <= 12'hb27;
      20'h09255: out <= 12'hb27;
      20'h09256: out <= 12'hf87;
      20'h09257: out <= 12'hb27;
      20'h09258: out <= 12'h000;
      20'h09259: out <= 12'h000;
      20'h0925a: out <= 12'h000;
      20'h0925b: out <= 12'h000;
      20'h0925c: out <= 12'h000;
      20'h0925d: out <= 12'h000;
      20'h0925e: out <= 12'h000;
      20'h0925f: out <= 12'h000;
      20'h09260: out <= 12'h8d0;
      20'h09261: out <= 12'h8d0;
      20'h09262: out <= 12'h000;
      20'h09263: out <= 12'h000;
      20'h09264: out <= 12'h000;
      20'h09265: out <= 12'h000;
      20'h09266: out <= 12'h000;
      20'h09267: out <= 12'h000;
      20'h09268: out <= 12'h8d0;
      20'h09269: out <= 12'h8d0;
      20'h0926a: out <= 12'h000;
      20'h0926b: out <= 12'h000;
      20'h0926c: out <= 12'h000;
      20'h0926d: out <= 12'h000;
      20'h0926e: out <= 12'h000;
      20'h0926f: out <= 12'h8d0;
      20'h09270: out <= 12'h8d0;
      20'h09271: out <= 12'h000;
      20'h09272: out <= 12'h000;
      20'h09273: out <= 12'h000;
      20'h09274: out <= 12'h000;
      20'h09275: out <= 12'h8d0;
      20'h09276: out <= 12'h8d0;
      20'h09277: out <= 12'h000;
      20'h09278: out <= 12'h000;
      20'h09279: out <= 12'h8d0;
      20'h0927a: out <= 12'h8d0;
      20'h0927b: out <= 12'h000;
      20'h0927c: out <= 12'h000;
      20'h0927d: out <= 12'h000;
      20'h0927e: out <= 12'h8d0;
      20'h0927f: out <= 12'h8d0;
      20'h09280: out <= 12'h8d0;
      20'h09281: out <= 12'h000;
      20'h09282: out <= 12'h000;
      20'h09283: out <= 12'h000;
      20'h09284: out <= 12'h000;
      20'h09285: out <= 12'h000;
      20'h09286: out <= 12'h000;
      20'h09287: out <= 12'h000;
      20'h09288: out <= 12'h000;
      20'h09289: out <= 12'h000;
      20'h0928a: out <= 12'h000;
      20'h0928b: out <= 12'h000;
      20'h0928c: out <= 12'h000;
      20'h0928d: out <= 12'h000;
      20'h0928e: out <= 12'h000;
      20'h0928f: out <= 12'h000;
      20'h09290: out <= 12'h222;
      20'h09291: out <= 12'h666;
      20'h09292: out <= 12'hbbb;
      20'h09293: out <= 12'h666;
      20'h09294: out <= 12'hfff;
      20'h09295: out <= 12'hbbb;
      20'h09296: out <= 12'hbbb;
      20'h09297: out <= 12'hbbb;
      20'h09298: out <= 12'h666;
      20'h09299: out <= 12'h666;
      20'h0929a: out <= 12'h666;
      20'h0929b: out <= 12'hbbb;
      20'h0929c: out <= 12'hbbb;
      20'h0929d: out <= 12'hbbb;
      20'h0929e: out <= 12'hbbb;
      20'h0929f: out <= 12'hbbb;
      20'h092a0: out <= 12'h000;
      20'h092a1: out <= 12'h666;
      20'h092a2: out <= 12'hbbb;
      20'h092a3: out <= 12'h666;
      20'h092a4: out <= 12'hbbb;
      20'h092a5: out <= 12'hbbb;
      20'h092a6: out <= 12'hbbb;
      20'h092a7: out <= 12'h666;
      20'h092a8: out <= 12'h666;
      20'h092a9: out <= 12'h666;
      20'h092aa: out <= 12'h666;
      20'h092ab: out <= 12'hbbb;
      20'h092ac: out <= 12'hbbb;
      20'h092ad: out <= 12'hbbb;
      20'h092ae: out <= 12'hbbb;
      20'h092af: out <= 12'hbbb;
      20'h092b0: out <= 12'h222;
      20'h092b1: out <= 12'h666;
      20'h092b2: out <= 12'hfff;
      20'h092b3: out <= 12'h666;
      20'h092b4: out <= 12'hbbb;
      20'h092b5: out <= 12'hbbb;
      20'h092b6: out <= 12'h666;
      20'h092b7: out <= 12'h666;
      20'h092b8: out <= 12'h666;
      20'h092b9: out <= 12'hbbb;
      20'h092ba: out <= 12'h666;
      20'h092bb: out <= 12'hbbb;
      20'h092bc: out <= 12'hbbb;
      20'h092bd: out <= 12'h666;
      20'h092be: out <= 12'hfff;
      20'h092bf: out <= 12'h666;
      20'h092c0: out <= 12'h000;
      20'h092c1: out <= 12'h666;
      20'h092c2: out <= 12'h666;
      20'h092c3: out <= 12'h666;
      20'h092c4: out <= 12'hbbb;
      20'h092c5: out <= 12'hbbb;
      20'h092c6: out <= 12'h666;
      20'h092c7: out <= 12'h666;
      20'h092c8: out <= 12'h666;
      20'h092c9: out <= 12'h666;
      20'h092ca: out <= 12'h666;
      20'h092cb: out <= 12'hbbb;
      20'h092cc: out <= 12'hbbb;
      20'h092cd: out <= 12'h666;
      20'h092ce: out <= 12'h666;
      20'h092cf: out <= 12'h666;
      20'h092d0: out <= 12'hbbb;
      20'h092d1: out <= 12'hbbb;
      20'h092d2: out <= 12'hbbb;
      20'h092d3: out <= 12'hbbb;
      20'h092d4: out <= 12'hbbb;
      20'h092d5: out <= 12'h666;
      20'h092d6: out <= 12'h666;
      20'h092d7: out <= 12'h666;
      20'h092d8: out <= 12'hbbb;
      20'h092d9: out <= 12'hbbb;
      20'h092da: out <= 12'hbbb;
      20'h092db: out <= 12'hfff;
      20'h092dc: out <= 12'h666;
      20'h092dd: out <= 12'hbbb;
      20'h092de: out <= 12'h666;
      20'h092df: out <= 12'h222;
      20'h092e0: out <= 12'hbbb;
      20'h092e1: out <= 12'hbbb;
      20'h092e2: out <= 12'hbbb;
      20'h092e3: out <= 12'hbbb;
      20'h092e4: out <= 12'hbbb;
      20'h092e5: out <= 12'h666;
      20'h092e6: out <= 12'h666;
      20'h092e7: out <= 12'h666;
      20'h092e8: out <= 12'h666;
      20'h092e9: out <= 12'hbbb;
      20'h092ea: out <= 12'hbbb;
      20'h092eb: out <= 12'hbbb;
      20'h092ec: out <= 12'h666;
      20'h092ed: out <= 12'hbbb;
      20'h092ee: out <= 12'h666;
      20'h092ef: out <= 12'h000;
      20'h092f0: out <= 12'h222;
      20'h092f1: out <= 12'h666;
      20'h092f2: out <= 12'h666;
      20'h092f3: out <= 12'h666;
      20'h092f4: out <= 12'hbbb;
      20'h092f5: out <= 12'h666;
      20'h092f6: out <= 12'h666;
      20'h092f7: out <= 12'hbbb;
      20'h092f8: out <= 12'hbbb;
      20'h092f9: out <= 12'hfff;
      20'h092fa: out <= 12'h666;
      20'h092fb: out <= 12'h666;
      20'h092fc: out <= 12'hbbb;
      20'h092fd: out <= 12'h666;
      20'h092fe: out <= 12'h666;
      20'h092ff: out <= 12'h666;
      20'h09300: out <= 12'h000;
      20'h09301: out <= 12'h666;
      20'h09302: out <= 12'hfff;
      20'h09303: out <= 12'h666;
      20'h09304: out <= 12'hbbb;
      20'h09305: out <= 12'h666;
      20'h09306: out <= 12'h666;
      20'h09307: out <= 12'hbbb;
      20'h09308: out <= 12'hbbb;
      20'h09309: out <= 12'hbbb;
      20'h0930a: out <= 12'h666;
      20'h0930b: out <= 12'h666;
      20'h0930c: out <= 12'hbbb;
      20'h0930d: out <= 12'h666;
      20'h0930e: out <= 12'hfff;
      20'h0930f: out <= 12'h666;
      20'h09310: out <= 12'h603;
      20'h09311: out <= 12'h603;
      20'h09312: out <= 12'h603;
      20'h09313: out <= 12'h603;
      20'h09314: out <= 12'h603;
      20'h09315: out <= 12'h603;
      20'h09316: out <= 12'h603;
      20'h09317: out <= 12'h603;
      20'h09318: out <= 12'h603;
      20'h09319: out <= 12'h603;
      20'h0931a: out <= 12'h603;
      20'h0931b: out <= 12'h603;
      20'h0931c: out <= 12'h603;
      20'h0931d: out <= 12'h603;
      20'h0931e: out <= 12'h603;
      20'h0931f: out <= 12'h603;
      20'h09320: out <= 12'h603;
      20'h09321: out <= 12'h603;
      20'h09322: out <= 12'h603;
      20'h09323: out <= 12'h603;
      20'h09324: out <= 12'h603;
      20'h09325: out <= 12'h603;
      20'h09326: out <= 12'h603;
      20'h09327: out <= 12'h603;
      20'h09328: out <= 12'h603;
      20'h09329: out <= 12'h603;
      20'h0932a: out <= 12'h603;
      20'h0932b: out <= 12'h603;
      20'h0932c: out <= 12'h603;
      20'h0932d: out <= 12'h603;
      20'h0932e: out <= 12'h603;
      20'h0932f: out <= 12'h603;
      20'h09330: out <= 12'h603;
      20'h09331: out <= 12'h603;
      20'h09332: out <= 12'h603;
      20'h09333: out <= 12'h603;
      20'h09334: out <= 12'h603;
      20'h09335: out <= 12'h603;
      20'h09336: out <= 12'h603;
      20'h09337: out <= 12'h603;
      20'h09338: out <= 12'h603;
      20'h09339: out <= 12'h603;
      20'h0933a: out <= 12'h603;
      20'h0933b: out <= 12'h603;
      20'h0933c: out <= 12'h603;
      20'h0933d: out <= 12'h603;
      20'h0933e: out <= 12'h603;
      20'h0933f: out <= 12'h603;
      20'h09340: out <= 12'h603;
      20'h09341: out <= 12'h603;
      20'h09342: out <= 12'h603;
      20'h09343: out <= 12'h603;
      20'h09344: out <= 12'h603;
      20'h09345: out <= 12'h603;
      20'h09346: out <= 12'h603;
      20'h09347: out <= 12'h603;
      20'h09348: out <= 12'h603;
      20'h09349: out <= 12'h603;
      20'h0934a: out <= 12'h603;
      20'h0934b: out <= 12'h603;
      20'h0934c: out <= 12'h603;
      20'h0934d: out <= 12'h603;
      20'h0934e: out <= 12'h603;
      20'h0934f: out <= 12'h603;
      20'h09350: out <= 12'h603;
      20'h09351: out <= 12'h603;
      20'h09352: out <= 12'h603;
      20'h09353: out <= 12'h603;
      20'h09354: out <= 12'h603;
      20'h09355: out <= 12'h603;
      20'h09356: out <= 12'h603;
      20'h09357: out <= 12'h603;
      20'h09358: out <= 12'h603;
      20'h09359: out <= 12'h603;
      20'h0935a: out <= 12'h603;
      20'h0935b: out <= 12'h603;
      20'h0935c: out <= 12'h603;
      20'h0935d: out <= 12'h603;
      20'h0935e: out <= 12'h603;
      20'h0935f: out <= 12'h603;
      20'h09360: out <= 12'h603;
      20'h09361: out <= 12'h603;
      20'h09362: out <= 12'h603;
      20'h09363: out <= 12'h603;
      20'h09364: out <= 12'h603;
      20'h09365: out <= 12'h603;
      20'h09366: out <= 12'h603;
      20'h09367: out <= 12'h603;
      20'h09368: out <= 12'hee9;
      20'h09369: out <= 12'hf87;
      20'h0936a: out <= 12'hf87;
      20'h0936b: out <= 12'hf87;
      20'h0936c: out <= 12'hf87;
      20'h0936d: out <= 12'hf87;
      20'h0936e: out <= 12'hf87;
      20'h0936f: out <= 12'hb27;
      20'h09370: out <= 12'h000;
      20'h09371: out <= 12'h000;
      20'h09372: out <= 12'h000;
      20'h09373: out <= 12'h000;
      20'h09374: out <= 12'h000;
      20'h09375: out <= 12'h000;
      20'h09376: out <= 12'h000;
      20'h09377: out <= 12'h000;
      20'h09378: out <= 12'h8d0;
      20'h09379: out <= 12'h8d0;
      20'h0937a: out <= 12'h8d0;
      20'h0937b: out <= 12'h8d0;
      20'h0937c: out <= 12'h8d0;
      20'h0937d: out <= 12'h8d0;
      20'h0937e: out <= 12'h8d0;
      20'h0937f: out <= 12'h000;
      20'h09380: out <= 12'h8d0;
      20'h09381: out <= 12'h8d0;
      20'h09382: out <= 12'h000;
      20'h09383: out <= 12'h000;
      20'h09384: out <= 12'h000;
      20'h09385: out <= 12'h000;
      20'h09386: out <= 12'h000;
      20'h09387: out <= 12'h8d0;
      20'h09388: out <= 12'h8d0;
      20'h09389: out <= 12'h8d0;
      20'h0938a: out <= 12'h8d0;
      20'h0938b: out <= 12'h8d0;
      20'h0938c: out <= 12'h000;
      20'h0938d: out <= 12'h8d0;
      20'h0938e: out <= 12'h8d0;
      20'h0938f: out <= 12'h000;
      20'h09390: out <= 12'h000;
      20'h09391: out <= 12'h8d0;
      20'h09392: out <= 12'h8d0;
      20'h09393: out <= 12'h000;
      20'h09394: out <= 12'h000;
      20'h09395: out <= 12'h000;
      20'h09396: out <= 12'h8d0;
      20'h09397: out <= 12'h8d0;
      20'h09398: out <= 12'h8d0;
      20'h09399: out <= 12'h000;
      20'h0939a: out <= 12'h000;
      20'h0939b: out <= 12'h000;
      20'h0939c: out <= 12'h000;
      20'h0939d: out <= 12'h000;
      20'h0939e: out <= 12'h000;
      20'h0939f: out <= 12'h000;
      20'h093a0: out <= 12'h000;
      20'h093a1: out <= 12'h000;
      20'h093a2: out <= 12'h000;
      20'h093a3: out <= 12'h000;
      20'h093a4: out <= 12'h000;
      20'h093a5: out <= 12'h000;
      20'h093a6: out <= 12'h000;
      20'h093a7: out <= 12'h000;
      20'h093a8: out <= 12'h222;
      20'h093a9: out <= 12'h666;
      20'h093aa: out <= 12'h666;
      20'h093ab: out <= 12'h666;
      20'h093ac: out <= 12'hfff;
      20'h093ad: out <= 12'hfff;
      20'h093ae: out <= 12'hbbb;
      20'h093af: out <= 12'hbbb;
      20'h093b0: out <= 12'hbbb;
      20'h093b1: out <= 12'h666;
      20'h093b2: out <= 12'h666;
      20'h093b3: out <= 12'hfff;
      20'h093b4: out <= 12'hfff;
      20'h093b5: out <= 12'hfff;
      20'h093b6: out <= 12'hfff;
      20'h093b7: out <= 12'hfff;
      20'h093b8: out <= 12'h000;
      20'h093b9: out <= 12'h666;
      20'h093ba: out <= 12'h666;
      20'h093bb: out <= 12'h666;
      20'h093bc: out <= 12'hfff;
      20'h093bd: out <= 12'hbbb;
      20'h093be: out <= 12'hbbb;
      20'h093bf: out <= 12'hbbb;
      20'h093c0: out <= 12'h666;
      20'h093c1: out <= 12'h666;
      20'h093c2: out <= 12'h666;
      20'h093c3: out <= 12'hfff;
      20'h093c4: out <= 12'hfff;
      20'h093c5: out <= 12'hfff;
      20'h093c6: out <= 12'hfff;
      20'h093c7: out <= 12'hfff;
      20'h093c8: out <= 12'h222;
      20'h093c9: out <= 12'h666;
      20'h093ca: out <= 12'h666;
      20'h093cb: out <= 12'h666;
      20'h093cc: out <= 12'hbbb;
      20'h093cd: out <= 12'h666;
      20'h093ce: out <= 12'h666;
      20'h093cf: out <= 12'h666;
      20'h093d0: out <= 12'hbbb;
      20'h093d1: out <= 12'hbbb;
      20'h093d2: out <= 12'h666;
      20'h093d3: out <= 12'h666;
      20'h093d4: out <= 12'hbbb;
      20'h093d5: out <= 12'h666;
      20'h093d6: out <= 12'h666;
      20'h093d7: out <= 12'h666;
      20'h093d8: out <= 12'h000;
      20'h093d9: out <= 12'h666;
      20'h093da: out <= 12'hfff;
      20'h093db: out <= 12'h666;
      20'h093dc: out <= 12'hbbb;
      20'h093dd: out <= 12'h666;
      20'h093de: out <= 12'h666;
      20'h093df: out <= 12'h666;
      20'h093e0: out <= 12'h666;
      20'h093e1: out <= 12'hbbb;
      20'h093e2: out <= 12'h666;
      20'h093e3: out <= 12'h666;
      20'h093e4: out <= 12'hbbb;
      20'h093e5: out <= 12'h666;
      20'h093e6: out <= 12'hfff;
      20'h093e7: out <= 12'h666;
      20'h093e8: out <= 12'hfff;
      20'h093e9: out <= 12'hfff;
      20'h093ea: out <= 12'hfff;
      20'h093eb: out <= 12'hfff;
      20'h093ec: out <= 12'hfff;
      20'h093ed: out <= 12'h666;
      20'h093ee: out <= 12'h666;
      20'h093ef: out <= 12'hbbb;
      20'h093f0: out <= 12'hbbb;
      20'h093f1: out <= 12'hbbb;
      20'h093f2: out <= 12'hfff;
      20'h093f3: out <= 12'hfff;
      20'h093f4: out <= 12'h666;
      20'h093f5: out <= 12'h666;
      20'h093f6: out <= 12'h666;
      20'h093f7: out <= 12'h222;
      20'h093f8: out <= 12'hfff;
      20'h093f9: out <= 12'hfff;
      20'h093fa: out <= 12'hfff;
      20'h093fb: out <= 12'hfff;
      20'h093fc: out <= 12'hfff;
      20'h093fd: out <= 12'h666;
      20'h093fe: out <= 12'h666;
      20'h093ff: out <= 12'h666;
      20'h09400: out <= 12'hbbb;
      20'h09401: out <= 12'hbbb;
      20'h09402: out <= 12'hbbb;
      20'h09403: out <= 12'hfff;
      20'h09404: out <= 12'h666;
      20'h09405: out <= 12'h666;
      20'h09406: out <= 12'h666;
      20'h09407: out <= 12'h000;
      20'h09408: out <= 12'h222;
      20'h09409: out <= 12'h666;
      20'h0940a: out <= 12'hfff;
      20'h0940b: out <= 12'h666;
      20'h0940c: out <= 12'hbbb;
      20'h0940d: out <= 12'hbbb;
      20'h0940e: out <= 12'h666;
      20'h0940f: out <= 12'hbbb;
      20'h09410: out <= 12'hbbb;
      20'h09411: out <= 12'hbbb;
      20'h09412: out <= 12'h666;
      20'h09413: out <= 12'hbbb;
      20'h09414: out <= 12'hbbb;
      20'h09415: out <= 12'h666;
      20'h09416: out <= 12'hfff;
      20'h09417: out <= 12'h666;
      20'h09418: out <= 12'h000;
      20'h09419: out <= 12'h666;
      20'h0941a: out <= 12'h666;
      20'h0941b: out <= 12'h666;
      20'h0941c: out <= 12'hbbb;
      20'h0941d: out <= 12'hbbb;
      20'h0941e: out <= 12'h666;
      20'h0941f: out <= 12'h666;
      20'h09420: out <= 12'hbbb;
      20'h09421: out <= 12'hbbb;
      20'h09422: out <= 12'h666;
      20'h09423: out <= 12'hbbb;
      20'h09424: out <= 12'hbbb;
      20'h09425: out <= 12'h666;
      20'h09426: out <= 12'h666;
      20'h09427: out <= 12'h666;
      20'h09428: out <= 12'h603;
      20'h09429: out <= 12'h603;
      20'h0942a: out <= 12'h603;
      20'h0942b: out <= 12'h603;
      20'h0942c: out <= 12'h603;
      20'h0942d: out <= 12'h603;
      20'h0942e: out <= 12'h603;
      20'h0942f: out <= 12'h603;
      20'h09430: out <= 12'h603;
      20'h09431: out <= 12'h603;
      20'h09432: out <= 12'h603;
      20'h09433: out <= 12'h603;
      20'h09434: out <= 12'h603;
      20'h09435: out <= 12'h603;
      20'h09436: out <= 12'h603;
      20'h09437: out <= 12'h603;
      20'h09438: out <= 12'h603;
      20'h09439: out <= 12'h603;
      20'h0943a: out <= 12'h603;
      20'h0943b: out <= 12'h603;
      20'h0943c: out <= 12'h603;
      20'h0943d: out <= 12'h603;
      20'h0943e: out <= 12'h603;
      20'h0943f: out <= 12'h603;
      20'h09440: out <= 12'h603;
      20'h09441: out <= 12'h603;
      20'h09442: out <= 12'h603;
      20'h09443: out <= 12'h603;
      20'h09444: out <= 12'h603;
      20'h09445: out <= 12'h603;
      20'h09446: out <= 12'h603;
      20'h09447: out <= 12'h603;
      20'h09448: out <= 12'h603;
      20'h09449: out <= 12'h603;
      20'h0944a: out <= 12'h603;
      20'h0944b: out <= 12'h603;
      20'h0944c: out <= 12'h603;
      20'h0944d: out <= 12'h603;
      20'h0944e: out <= 12'h603;
      20'h0944f: out <= 12'h603;
      20'h09450: out <= 12'h603;
      20'h09451: out <= 12'h603;
      20'h09452: out <= 12'h603;
      20'h09453: out <= 12'h603;
      20'h09454: out <= 12'h603;
      20'h09455: out <= 12'h603;
      20'h09456: out <= 12'h603;
      20'h09457: out <= 12'h603;
      20'h09458: out <= 12'h603;
      20'h09459: out <= 12'h603;
      20'h0945a: out <= 12'h603;
      20'h0945b: out <= 12'h603;
      20'h0945c: out <= 12'h603;
      20'h0945d: out <= 12'h603;
      20'h0945e: out <= 12'h603;
      20'h0945f: out <= 12'h603;
      20'h09460: out <= 12'h603;
      20'h09461: out <= 12'h603;
      20'h09462: out <= 12'h603;
      20'h09463: out <= 12'h603;
      20'h09464: out <= 12'h603;
      20'h09465: out <= 12'h603;
      20'h09466: out <= 12'h603;
      20'h09467: out <= 12'h603;
      20'h09468: out <= 12'h603;
      20'h09469: out <= 12'h603;
      20'h0946a: out <= 12'h603;
      20'h0946b: out <= 12'h603;
      20'h0946c: out <= 12'h603;
      20'h0946d: out <= 12'h603;
      20'h0946e: out <= 12'h603;
      20'h0946f: out <= 12'h603;
      20'h09470: out <= 12'h603;
      20'h09471: out <= 12'h603;
      20'h09472: out <= 12'h603;
      20'h09473: out <= 12'h603;
      20'h09474: out <= 12'h603;
      20'h09475: out <= 12'h603;
      20'h09476: out <= 12'h603;
      20'h09477: out <= 12'h603;
      20'h09478: out <= 12'h603;
      20'h09479: out <= 12'h603;
      20'h0947a: out <= 12'h603;
      20'h0947b: out <= 12'h603;
      20'h0947c: out <= 12'h603;
      20'h0947d: out <= 12'h603;
      20'h0947e: out <= 12'h603;
      20'h0947f: out <= 12'h603;
      20'h09480: out <= 12'hb27;
      20'h09481: out <= 12'hb27;
      20'h09482: out <= 12'hb27;
      20'h09483: out <= 12'hb27;
      20'h09484: out <= 12'hb27;
      20'h09485: out <= 12'hb27;
      20'h09486: out <= 12'hb27;
      20'h09487: out <= 12'hb27;
      20'h09488: out <= 12'h000;
      20'h09489: out <= 12'h000;
      20'h0948a: out <= 12'h000;
      20'h0948b: out <= 12'h000;
      20'h0948c: out <= 12'h000;
      20'h0948d: out <= 12'h000;
      20'h0948e: out <= 12'h000;
      20'h0948f: out <= 12'h000;
      20'h09490: out <= 12'h000;
      20'h09491: out <= 12'h000;
      20'h09492: out <= 12'h000;
      20'h09493: out <= 12'h000;
      20'h09494: out <= 12'h000;
      20'h09495: out <= 12'h000;
      20'h09496: out <= 12'h000;
      20'h09497: out <= 12'h000;
      20'h09498: out <= 12'h000;
      20'h09499: out <= 12'h000;
      20'h0949a: out <= 12'h000;
      20'h0949b: out <= 12'h000;
      20'h0949c: out <= 12'h000;
      20'h0949d: out <= 12'h000;
      20'h0949e: out <= 12'h000;
      20'h0949f: out <= 12'h000;
      20'h094a0: out <= 12'h000;
      20'h094a1: out <= 12'h000;
      20'h094a2: out <= 12'h000;
      20'h094a3: out <= 12'h000;
      20'h094a4: out <= 12'h000;
      20'h094a5: out <= 12'h000;
      20'h094a6: out <= 12'h000;
      20'h094a7: out <= 12'h000;
      20'h094a8: out <= 12'h000;
      20'h094a9: out <= 12'h000;
      20'h094aa: out <= 12'h000;
      20'h094ab: out <= 12'h000;
      20'h094ac: out <= 12'h000;
      20'h094ad: out <= 12'h000;
      20'h094ae: out <= 12'h000;
      20'h094af: out <= 12'h000;
      20'h094b0: out <= 12'h000;
      20'h094b1: out <= 12'h000;
      20'h094b2: out <= 12'h000;
      20'h094b3: out <= 12'h000;
      20'h094b4: out <= 12'h000;
      20'h094b5: out <= 12'h000;
      20'h094b6: out <= 12'h000;
      20'h094b7: out <= 12'h000;
      20'h094b8: out <= 12'h000;
      20'h094b9: out <= 12'h000;
      20'h094ba: out <= 12'h000;
      20'h094bb: out <= 12'h000;
      20'h094bc: out <= 12'h000;
      20'h094bd: out <= 12'h000;
      20'h094be: out <= 12'h000;
      20'h094bf: out <= 12'h000;
      20'h094c0: out <= 12'h222;
      20'h094c1: out <= 12'h666;
      20'h094c2: out <= 12'hbbb;
      20'h094c3: out <= 12'h666;
      20'h094c4: out <= 12'hfff;
      20'h094c5: out <= 12'hfff;
      20'h094c6: out <= 12'hfff;
      20'h094c7: out <= 12'hbbb;
      20'h094c8: out <= 12'hbbb;
      20'h094c9: out <= 12'hbbb;
      20'h094ca: out <= 12'h666;
      20'h094cb: out <= 12'hbbb;
      20'h094cc: out <= 12'hbbb;
      20'h094cd: out <= 12'hbbb;
      20'h094ce: out <= 12'hbbb;
      20'h094cf: out <= 12'hbbb;
      20'h094d0: out <= 12'h000;
      20'h094d1: out <= 12'h666;
      20'h094d2: out <= 12'hbbb;
      20'h094d3: out <= 12'h666;
      20'h094d4: out <= 12'hfff;
      20'h094d5: out <= 12'hfff;
      20'h094d6: out <= 12'hbbb;
      20'h094d7: out <= 12'hbbb;
      20'h094d8: out <= 12'hbbb;
      20'h094d9: out <= 12'h666;
      20'h094da: out <= 12'h666;
      20'h094db: out <= 12'hbbb;
      20'h094dc: out <= 12'hbbb;
      20'h094dd: out <= 12'hbbb;
      20'h094de: out <= 12'hbbb;
      20'h094df: out <= 12'hbbb;
      20'h094e0: out <= 12'h222;
      20'h094e1: out <= 12'h666;
      20'h094e2: out <= 12'hfff;
      20'h094e3: out <= 12'h666;
      20'h094e4: out <= 12'hbbb;
      20'h094e5: out <= 12'hbbb;
      20'h094e6: out <= 12'h666;
      20'h094e7: out <= 12'hbbb;
      20'h094e8: out <= 12'hbbb;
      20'h094e9: out <= 12'hbbb;
      20'h094ea: out <= 12'h666;
      20'h094eb: out <= 12'hbbb;
      20'h094ec: out <= 12'hbbb;
      20'h094ed: out <= 12'h666;
      20'h094ee: out <= 12'hfff;
      20'h094ef: out <= 12'h666;
      20'h094f0: out <= 12'h000;
      20'h094f1: out <= 12'h666;
      20'h094f2: out <= 12'h666;
      20'h094f3: out <= 12'h666;
      20'h094f4: out <= 12'hbbb;
      20'h094f5: out <= 12'hbbb;
      20'h094f6: out <= 12'h666;
      20'h094f7: out <= 12'h666;
      20'h094f8: out <= 12'hbbb;
      20'h094f9: out <= 12'hbbb;
      20'h094fa: out <= 12'h666;
      20'h094fb: out <= 12'hbbb;
      20'h094fc: out <= 12'hbbb;
      20'h094fd: out <= 12'h666;
      20'h094fe: out <= 12'h666;
      20'h094ff: out <= 12'h666;
      20'h09500: out <= 12'hbbb;
      20'h09501: out <= 12'hbbb;
      20'h09502: out <= 12'hbbb;
      20'h09503: out <= 12'hbbb;
      20'h09504: out <= 12'hbbb;
      20'h09505: out <= 12'h666;
      20'h09506: out <= 12'hbbb;
      20'h09507: out <= 12'hbbb;
      20'h09508: out <= 12'hbbb;
      20'h09509: out <= 12'hfff;
      20'h0950a: out <= 12'hfff;
      20'h0950b: out <= 12'hfff;
      20'h0950c: out <= 12'h666;
      20'h0950d: out <= 12'hbbb;
      20'h0950e: out <= 12'h666;
      20'h0950f: out <= 12'h222;
      20'h09510: out <= 12'hbbb;
      20'h09511: out <= 12'hbbb;
      20'h09512: out <= 12'hbbb;
      20'h09513: out <= 12'hbbb;
      20'h09514: out <= 12'hbbb;
      20'h09515: out <= 12'h666;
      20'h09516: out <= 12'h666;
      20'h09517: out <= 12'hbbb;
      20'h09518: out <= 12'hbbb;
      20'h09519: out <= 12'hbbb;
      20'h0951a: out <= 12'hfff;
      20'h0951b: out <= 12'hfff;
      20'h0951c: out <= 12'h666;
      20'h0951d: out <= 12'hbbb;
      20'h0951e: out <= 12'h666;
      20'h0951f: out <= 12'h000;
      20'h09520: out <= 12'h222;
      20'h09521: out <= 12'h666;
      20'h09522: out <= 12'h666;
      20'h09523: out <= 12'h666;
      20'h09524: out <= 12'hbbb;
      20'h09525: out <= 12'h666;
      20'h09526: out <= 12'h666;
      20'h09527: out <= 12'h666;
      20'h09528: out <= 12'hbbb;
      20'h09529: out <= 12'hbbb;
      20'h0952a: out <= 12'h666;
      20'h0952b: out <= 12'h666;
      20'h0952c: out <= 12'hbbb;
      20'h0952d: out <= 12'h666;
      20'h0952e: out <= 12'h666;
      20'h0952f: out <= 12'h666;
      20'h09530: out <= 12'h000;
      20'h09531: out <= 12'h666;
      20'h09532: out <= 12'hfff;
      20'h09533: out <= 12'h666;
      20'h09534: out <= 12'hbbb;
      20'h09535: out <= 12'h666;
      20'h09536: out <= 12'h666;
      20'h09537: out <= 12'h666;
      20'h09538: out <= 12'h666;
      20'h09539: out <= 12'hbbb;
      20'h0953a: out <= 12'h666;
      20'h0953b: out <= 12'h666;
      20'h0953c: out <= 12'hbbb;
      20'h0953d: out <= 12'h666;
      20'h0953e: out <= 12'hfff;
      20'h0953f: out <= 12'h666;
      20'h09540: out <= 12'h603;
      20'h09541: out <= 12'h603;
      20'h09542: out <= 12'h603;
      20'h09543: out <= 12'h603;
      20'h09544: out <= 12'h000;
      20'h09545: out <= 12'hf87;
      20'h09546: out <= 12'hf87;
      20'h09547: out <= 12'hf87;
      20'h09548: out <= 12'hf87;
      20'h09549: out <= 12'hf87;
      20'h0954a: out <= 12'h000;
      20'h0954b: out <= 12'h000;
      20'h0954c: out <= 12'h000;
      20'h0954d: out <= 12'h000;
      20'h0954e: out <= 12'h000;
      20'h0954f: out <= 12'hf87;
      20'h09550: out <= 12'hf87;
      20'h09551: out <= 12'h000;
      20'h09552: out <= 12'h000;
      20'h09553: out <= 12'h000;
      20'h09554: out <= 12'h000;
      20'h09555: out <= 12'hf87;
      20'h09556: out <= 12'hf87;
      20'h09557: out <= 12'hf87;
      20'h09558: out <= 12'hf87;
      20'h09559: out <= 12'hf87;
      20'h0955a: out <= 12'h000;
      20'h0955b: out <= 12'h000;
      20'h0955c: out <= 12'h000;
      20'h0955d: out <= 12'hf87;
      20'h0955e: out <= 12'hf87;
      20'h0955f: out <= 12'hf87;
      20'h09560: out <= 12'hf87;
      20'h09561: out <= 12'hf87;
      20'h09562: out <= 12'h000;
      20'h09563: out <= 12'h000;
      20'h09564: out <= 12'h000;
      20'h09565: out <= 12'h000;
      20'h09566: out <= 12'h000;
      20'h09567: out <= 12'hf87;
      20'h09568: out <= 12'hf87;
      20'h09569: out <= 12'hf87;
      20'h0956a: out <= 12'h000;
      20'h0956b: out <= 12'h000;
      20'h0956c: out <= 12'hf87;
      20'h0956d: out <= 12'hf87;
      20'h0956e: out <= 12'hf87;
      20'h0956f: out <= 12'hf87;
      20'h09570: out <= 12'hf87;
      20'h09571: out <= 12'hf87;
      20'h09572: out <= 12'hf87;
      20'h09573: out <= 12'h000;
      20'h09574: out <= 12'h000;
      20'h09575: out <= 12'h000;
      20'h09576: out <= 12'hf87;
      20'h09577: out <= 12'hf87;
      20'h09578: out <= 12'hf87;
      20'h09579: out <= 12'hf87;
      20'h0957a: out <= 12'h000;
      20'h0957b: out <= 12'h000;
      20'h0957c: out <= 12'hf87;
      20'h0957d: out <= 12'hf87;
      20'h0957e: out <= 12'hf87;
      20'h0957f: out <= 12'hf87;
      20'h09580: out <= 12'hf87;
      20'h09581: out <= 12'hf87;
      20'h09582: out <= 12'hf87;
      20'h09583: out <= 12'h000;
      20'h09584: out <= 12'h000;
      20'h09585: out <= 12'hf87;
      20'h09586: out <= 12'hf87;
      20'h09587: out <= 12'hf87;
      20'h09588: out <= 12'hf87;
      20'h09589: out <= 12'hf87;
      20'h0958a: out <= 12'h000;
      20'h0958b: out <= 12'h000;
      20'h0958c: out <= 12'h000;
      20'h0958d: out <= 12'hf87;
      20'h0958e: out <= 12'hf87;
      20'h0958f: out <= 12'hf87;
      20'h09590: out <= 12'hf87;
      20'h09591: out <= 12'hf87;
      20'h09592: out <= 12'h000;
      20'h09593: out <= 12'h000;
      20'h09594: out <= 12'h603;
      20'h09595: out <= 12'h603;
      20'h09596: out <= 12'h603;
      20'h09597: out <= 12'h603;
      20'h09598: out <= 12'hee9;
      20'h09599: out <= 12'hee9;
      20'h0959a: out <= 12'hee9;
      20'h0959b: out <= 12'hee9;
      20'h0959c: out <= 12'hee9;
      20'h0959d: out <= 12'hee9;
      20'h0959e: out <= 12'hee9;
      20'h0959f: out <= 12'hb27;
      20'h095a0: out <= 12'h000;
      20'h095a1: out <= 12'h000;
      20'h095a2: out <= 12'h000;
      20'h095a3: out <= 12'h000;
      20'h095a4: out <= 12'h000;
      20'h095a5: out <= 12'h000;
      20'h095a6: out <= 12'h000;
      20'h095a7: out <= 12'h000;
      20'h095a8: out <= 12'h000;
      20'h095a9: out <= 12'h000;
      20'h095aa: out <= 12'h000;
      20'h095ab: out <= 12'h000;
      20'h095ac: out <= 12'h000;
      20'h095ad: out <= 12'h000;
      20'h095ae: out <= 12'h000;
      20'h095af: out <= 12'hc7f;
      20'h095b0: out <= 12'hfff;
      20'h095b1: out <= 12'hc7f;
      20'h095b2: out <= 12'h000;
      20'h095b3: out <= 12'h000;
      20'h095b4: out <= 12'h000;
      20'h095b5: out <= 12'h000;
      20'h095b6: out <= 12'h000;
      20'h095b7: out <= 12'h000;
      20'h095b8: out <= 12'h000;
      20'h095b9: out <= 12'h000;
      20'h095ba: out <= 12'h000;
      20'h095bb: out <= 12'h000;
      20'h095bc: out <= 12'h000;
      20'h095bd: out <= 12'h000;
      20'h095be: out <= 12'h000;
      20'h095bf: out <= 12'h000;
      20'h095c0: out <= 12'h000;
      20'h095c1: out <= 12'h000;
      20'h095c2: out <= 12'h000;
      20'h095c3: out <= 12'h000;
      20'h095c4: out <= 12'h000;
      20'h095c5: out <= 12'h000;
      20'h095c6: out <= 12'h000;
      20'h095c7: out <= 12'h000;
      20'h095c8: out <= 12'h000;
      20'h095c9: out <= 12'h000;
      20'h095ca: out <= 12'h000;
      20'h095cb: out <= 12'h000;
      20'h095cc: out <= 12'h000;
      20'h095cd: out <= 12'h000;
      20'h095ce: out <= 12'h000;
      20'h095cf: out <= 12'h000;
      20'h095d0: out <= 12'h000;
      20'h095d1: out <= 12'h000;
      20'h095d2: out <= 12'h000;
      20'h095d3: out <= 12'h000;
      20'h095d4: out <= 12'h000;
      20'h095d5: out <= 12'h000;
      20'h095d6: out <= 12'h000;
      20'h095d7: out <= 12'h000;
      20'h095d8: out <= 12'h222;
      20'h095d9: out <= 12'h666;
      20'h095da: out <= 12'hfff;
      20'h095db: out <= 12'h666;
      20'h095dc: out <= 12'h666;
      20'h095dd: out <= 12'h666;
      20'h095de: out <= 12'h666;
      20'h095df: out <= 12'h666;
      20'h095e0: out <= 12'h666;
      20'h095e1: out <= 12'h666;
      20'h095e2: out <= 12'h666;
      20'h095e3: out <= 12'h666;
      20'h095e4: out <= 12'h666;
      20'h095e5: out <= 12'h222;
      20'h095e6: out <= 12'h222;
      20'h095e7: out <= 12'hbbb;
      20'h095e8: out <= 12'h000;
      20'h095e9: out <= 12'h666;
      20'h095ea: out <= 12'hfff;
      20'h095eb: out <= 12'h666;
      20'h095ec: out <= 12'h666;
      20'h095ed: out <= 12'h666;
      20'h095ee: out <= 12'h666;
      20'h095ef: out <= 12'h666;
      20'h095f0: out <= 12'h666;
      20'h095f1: out <= 12'h666;
      20'h095f2: out <= 12'h666;
      20'h095f3: out <= 12'h666;
      20'h095f4: out <= 12'h666;
      20'h095f5: out <= 12'h000;
      20'h095f6: out <= 12'h000;
      20'h095f7: out <= 12'hbbb;
      20'h095f8: out <= 12'h222;
      20'h095f9: out <= 12'h666;
      20'h095fa: out <= 12'h666;
      20'h095fb: out <= 12'h666;
      20'h095fc: out <= 12'hbbb;
      20'h095fd: out <= 12'h666;
      20'h095fe: out <= 12'h666;
      20'h095ff: out <= 12'hbbb;
      20'h09600: out <= 12'hbbb;
      20'h09601: out <= 12'hfff;
      20'h09602: out <= 12'h666;
      20'h09603: out <= 12'h666;
      20'h09604: out <= 12'hbbb;
      20'h09605: out <= 12'h666;
      20'h09606: out <= 12'h666;
      20'h09607: out <= 12'h666;
      20'h09608: out <= 12'h000;
      20'h09609: out <= 12'h666;
      20'h0960a: out <= 12'hfff;
      20'h0960b: out <= 12'h666;
      20'h0960c: out <= 12'hbbb;
      20'h0960d: out <= 12'h666;
      20'h0960e: out <= 12'h666;
      20'h0960f: out <= 12'hbbb;
      20'h09610: out <= 12'hbbb;
      20'h09611: out <= 12'hbbb;
      20'h09612: out <= 12'h666;
      20'h09613: out <= 12'h666;
      20'h09614: out <= 12'hbbb;
      20'h09615: out <= 12'h666;
      20'h09616: out <= 12'hfff;
      20'h09617: out <= 12'h666;
      20'h09618: out <= 12'hbbb;
      20'h09619: out <= 12'h222;
      20'h0961a: out <= 12'h222;
      20'h0961b: out <= 12'h666;
      20'h0961c: out <= 12'h666;
      20'h0961d: out <= 12'h666;
      20'h0961e: out <= 12'h666;
      20'h0961f: out <= 12'h666;
      20'h09620: out <= 12'h666;
      20'h09621: out <= 12'h666;
      20'h09622: out <= 12'h666;
      20'h09623: out <= 12'h666;
      20'h09624: out <= 12'h666;
      20'h09625: out <= 12'hfff;
      20'h09626: out <= 12'h666;
      20'h09627: out <= 12'h222;
      20'h09628: out <= 12'hbbb;
      20'h09629: out <= 12'h000;
      20'h0962a: out <= 12'h000;
      20'h0962b: out <= 12'h666;
      20'h0962c: out <= 12'h666;
      20'h0962d: out <= 12'h666;
      20'h0962e: out <= 12'h666;
      20'h0962f: out <= 12'h666;
      20'h09630: out <= 12'h666;
      20'h09631: out <= 12'h666;
      20'h09632: out <= 12'h666;
      20'h09633: out <= 12'h666;
      20'h09634: out <= 12'h666;
      20'h09635: out <= 12'hfff;
      20'h09636: out <= 12'h666;
      20'h09637: out <= 12'h000;
      20'h09638: out <= 12'h222;
      20'h09639: out <= 12'h666;
      20'h0963a: out <= 12'hfff;
      20'h0963b: out <= 12'h666;
      20'h0963c: out <= 12'hbbb;
      20'h0963d: out <= 12'hbbb;
      20'h0963e: out <= 12'h666;
      20'h0963f: out <= 12'h666;
      20'h09640: out <= 12'h666;
      20'h09641: out <= 12'hbbb;
      20'h09642: out <= 12'h666;
      20'h09643: out <= 12'hbbb;
      20'h09644: out <= 12'hbbb;
      20'h09645: out <= 12'h666;
      20'h09646: out <= 12'hfff;
      20'h09647: out <= 12'h666;
      20'h09648: out <= 12'h000;
      20'h09649: out <= 12'h666;
      20'h0964a: out <= 12'h666;
      20'h0964b: out <= 12'h666;
      20'h0964c: out <= 12'hbbb;
      20'h0964d: out <= 12'hbbb;
      20'h0964e: out <= 12'h666;
      20'h0964f: out <= 12'h666;
      20'h09650: out <= 12'h666;
      20'h09651: out <= 12'h666;
      20'h09652: out <= 12'h666;
      20'h09653: out <= 12'hbbb;
      20'h09654: out <= 12'hbbb;
      20'h09655: out <= 12'h666;
      20'h09656: out <= 12'h666;
      20'h09657: out <= 12'h666;
      20'h09658: out <= 12'h603;
      20'h09659: out <= 12'h603;
      20'h0965a: out <= 12'h603;
      20'h0965b: out <= 12'h603;
      20'h0965c: out <= 12'hf87;
      20'h0965d: out <= 12'hf87;
      20'h0965e: out <= 12'h000;
      20'h0965f: out <= 12'h000;
      20'h09660: out <= 12'h000;
      20'h09661: out <= 12'hf87;
      20'h09662: out <= 12'hf87;
      20'h09663: out <= 12'h000;
      20'h09664: out <= 12'h000;
      20'h09665: out <= 12'h000;
      20'h09666: out <= 12'hf87;
      20'h09667: out <= 12'hf87;
      20'h09668: out <= 12'hf87;
      20'h09669: out <= 12'h000;
      20'h0966a: out <= 12'h000;
      20'h0966b: out <= 12'h000;
      20'h0966c: out <= 12'hf87;
      20'h0966d: out <= 12'hf87;
      20'h0966e: out <= 12'h000;
      20'h0966f: out <= 12'h000;
      20'h09670: out <= 12'h000;
      20'h09671: out <= 12'hf87;
      20'h09672: out <= 12'hf87;
      20'h09673: out <= 12'h000;
      20'h09674: out <= 12'hf87;
      20'h09675: out <= 12'hf87;
      20'h09676: out <= 12'h000;
      20'h09677: out <= 12'h000;
      20'h09678: out <= 12'h000;
      20'h09679: out <= 12'hf87;
      20'h0967a: out <= 12'hf87;
      20'h0967b: out <= 12'h000;
      20'h0967c: out <= 12'h000;
      20'h0967d: out <= 12'h000;
      20'h0967e: out <= 12'hf87;
      20'h0967f: out <= 12'hf87;
      20'h09680: out <= 12'hf87;
      20'h09681: out <= 12'hf87;
      20'h09682: out <= 12'h000;
      20'h09683: out <= 12'h000;
      20'h09684: out <= 12'hf87;
      20'h09685: out <= 12'hf87;
      20'h09686: out <= 12'h000;
      20'h09687: out <= 12'h000;
      20'h09688: out <= 12'h000;
      20'h09689: out <= 12'h000;
      20'h0968a: out <= 12'h000;
      20'h0968b: out <= 12'h000;
      20'h0968c: out <= 12'h000;
      20'h0968d: out <= 12'hf87;
      20'h0968e: out <= 12'hf87;
      20'h0968f: out <= 12'h000;
      20'h09690: out <= 12'h000;
      20'h09691: out <= 12'h000;
      20'h09692: out <= 12'h000;
      20'h09693: out <= 12'h000;
      20'h09694: out <= 12'hf87;
      20'h09695: out <= 12'hf87;
      20'h09696: out <= 12'h000;
      20'h09697: out <= 12'h000;
      20'h09698: out <= 12'h000;
      20'h09699: out <= 12'hf87;
      20'h0969a: out <= 12'hf87;
      20'h0969b: out <= 12'h000;
      20'h0969c: out <= 12'hf87;
      20'h0969d: out <= 12'hf87;
      20'h0969e: out <= 12'h000;
      20'h0969f: out <= 12'h000;
      20'h096a0: out <= 12'h000;
      20'h096a1: out <= 12'hf87;
      20'h096a2: out <= 12'hf87;
      20'h096a3: out <= 12'h000;
      20'h096a4: out <= 12'hf87;
      20'h096a5: out <= 12'hf87;
      20'h096a6: out <= 12'h000;
      20'h096a7: out <= 12'h000;
      20'h096a8: out <= 12'h000;
      20'h096a9: out <= 12'hf87;
      20'h096aa: out <= 12'hf87;
      20'h096ab: out <= 12'h000;
      20'h096ac: out <= 12'h603;
      20'h096ad: out <= 12'h603;
      20'h096ae: out <= 12'h603;
      20'h096af: out <= 12'h603;
      20'h096b0: out <= 12'hee9;
      20'h096b1: out <= 12'hf87;
      20'h096b2: out <= 12'hf87;
      20'h096b3: out <= 12'hf87;
      20'h096b4: out <= 12'hf87;
      20'h096b5: out <= 12'hf87;
      20'h096b6: out <= 12'hf87;
      20'h096b7: out <= 12'hb27;
      20'h096b8: out <= 12'h000;
      20'h096b9: out <= 12'h000;
      20'h096ba: out <= 12'h000;
      20'h096bb: out <= 12'h000;
      20'h096bc: out <= 12'h000;
      20'h096bd: out <= 12'h000;
      20'h096be: out <= 12'h000;
      20'h096bf: out <= 12'h000;
      20'h096c0: out <= 12'h000;
      20'h096c1: out <= 12'h000;
      20'h096c2: out <= 12'h000;
      20'h096c3: out <= 12'h000;
      20'h096c4: out <= 12'h000;
      20'h096c5: out <= 12'h000;
      20'h096c6: out <= 12'h000;
      20'h096c7: out <= 12'h72f;
      20'h096c8: out <= 12'hfff;
      20'h096c9: out <= 12'h72f;
      20'h096ca: out <= 12'h000;
      20'h096cb: out <= 12'h000;
      20'h096cc: out <= 12'h000;
      20'h096cd: out <= 12'h000;
      20'h096ce: out <= 12'h000;
      20'h096cf: out <= 12'h000;
      20'h096d0: out <= 12'h000;
      20'h096d1: out <= 12'h000;
      20'h096d2: out <= 12'h000;
      20'h096d3: out <= 12'h000;
      20'h096d4: out <= 12'h000;
      20'h096d5: out <= 12'h000;
      20'h096d6: out <= 12'h000;
      20'h096d7: out <= 12'h000;
      20'h096d8: out <= 12'h000;
      20'h096d9: out <= 12'h000;
      20'h096da: out <= 12'h000;
      20'h096db: out <= 12'h000;
      20'h096dc: out <= 12'h000;
      20'h096dd: out <= 12'h000;
      20'h096de: out <= 12'h000;
      20'h096df: out <= 12'h000;
      20'h096e0: out <= 12'h000;
      20'h096e1: out <= 12'h000;
      20'h096e2: out <= 12'h000;
      20'h096e3: out <= 12'h000;
      20'h096e4: out <= 12'h000;
      20'h096e5: out <= 12'h000;
      20'h096e6: out <= 12'h000;
      20'h096e7: out <= 12'h000;
      20'h096e8: out <= 12'h000;
      20'h096e9: out <= 12'h000;
      20'h096ea: out <= 12'h000;
      20'h096eb: out <= 12'h000;
      20'h096ec: out <= 12'h000;
      20'h096ed: out <= 12'h000;
      20'h096ee: out <= 12'h000;
      20'h096ef: out <= 12'h000;
      20'h096f0: out <= 12'h222;
      20'h096f1: out <= 12'h222;
      20'h096f2: out <= 12'h666;
      20'h096f3: out <= 12'hfff;
      20'h096f4: out <= 12'hfff;
      20'h096f5: out <= 12'hbbb;
      20'h096f6: out <= 12'h666;
      20'h096f7: out <= 12'hbbb;
      20'h096f8: out <= 12'h666;
      20'h096f9: out <= 12'hbbb;
      20'h096fa: out <= 12'hfff;
      20'h096fb: out <= 12'hfff;
      20'h096fc: out <= 12'h666;
      20'h096fd: out <= 12'h222;
      20'h096fe: out <= 12'h222;
      20'h096ff: out <= 12'h222;
      20'h09700: out <= 12'h000;
      20'h09701: out <= 12'h000;
      20'h09702: out <= 12'h666;
      20'h09703: out <= 12'hfff;
      20'h09704: out <= 12'hfff;
      20'h09705: out <= 12'hbbb;
      20'h09706: out <= 12'h666;
      20'h09707: out <= 12'hbbb;
      20'h09708: out <= 12'h666;
      20'h09709: out <= 12'hbbb;
      20'h0970a: out <= 12'hfff;
      20'h0970b: out <= 12'hfff;
      20'h0970c: out <= 12'h666;
      20'h0970d: out <= 12'h000;
      20'h0970e: out <= 12'h000;
      20'h0970f: out <= 12'h000;
      20'h09710: out <= 12'h222;
      20'h09711: out <= 12'h666;
      20'h09712: out <= 12'hfff;
      20'h09713: out <= 12'h666;
      20'h09714: out <= 12'hbbb;
      20'h09715: out <= 12'hbbb;
      20'h09716: out <= 12'h666;
      20'h09717: out <= 12'hbbb;
      20'h09718: out <= 12'hfff;
      20'h09719: out <= 12'hfff;
      20'h0971a: out <= 12'h666;
      20'h0971b: out <= 12'hbbb;
      20'h0971c: out <= 12'hbbb;
      20'h0971d: out <= 12'h666;
      20'h0971e: out <= 12'hfff;
      20'h0971f: out <= 12'h666;
      20'h09720: out <= 12'h000;
      20'h09721: out <= 12'h666;
      20'h09722: out <= 12'h666;
      20'h09723: out <= 12'h666;
      20'h09724: out <= 12'hbbb;
      20'h09725: out <= 12'hbbb;
      20'h09726: out <= 12'h666;
      20'h09727: out <= 12'hbbb;
      20'h09728: out <= 12'hbbb;
      20'h09729: out <= 12'hfff;
      20'h0972a: out <= 12'h666;
      20'h0972b: out <= 12'hbbb;
      20'h0972c: out <= 12'hbbb;
      20'h0972d: out <= 12'h666;
      20'h0972e: out <= 12'h666;
      20'h0972f: out <= 12'h666;
      20'h09730: out <= 12'h222;
      20'h09731: out <= 12'h222;
      20'h09732: out <= 12'h222;
      20'h09733: out <= 12'h666;
      20'h09734: out <= 12'hfff;
      20'h09735: out <= 12'hfff;
      20'h09736: out <= 12'hbbb;
      20'h09737: out <= 12'h666;
      20'h09738: out <= 12'hbbb;
      20'h09739: out <= 12'h666;
      20'h0973a: out <= 12'hbbb;
      20'h0973b: out <= 12'hfff;
      20'h0973c: out <= 12'hfff;
      20'h0973d: out <= 12'h666;
      20'h0973e: out <= 12'h222;
      20'h0973f: out <= 12'h222;
      20'h09740: out <= 12'h000;
      20'h09741: out <= 12'h000;
      20'h09742: out <= 12'h000;
      20'h09743: out <= 12'h666;
      20'h09744: out <= 12'hfff;
      20'h09745: out <= 12'hfff;
      20'h09746: out <= 12'hbbb;
      20'h09747: out <= 12'h666;
      20'h09748: out <= 12'hbbb;
      20'h09749: out <= 12'h666;
      20'h0974a: out <= 12'hbbb;
      20'h0974b: out <= 12'hfff;
      20'h0974c: out <= 12'hfff;
      20'h0974d: out <= 12'h666;
      20'h0974e: out <= 12'h000;
      20'h0974f: out <= 12'h000;
      20'h09750: out <= 12'h222;
      20'h09751: out <= 12'h666;
      20'h09752: out <= 12'h666;
      20'h09753: out <= 12'h666;
      20'h09754: out <= 12'hbbb;
      20'h09755: out <= 12'hfff;
      20'h09756: out <= 12'h666;
      20'h09757: out <= 12'h666;
      20'h09758: out <= 12'h666;
      20'h09759: out <= 12'h666;
      20'h0975a: out <= 12'h666;
      20'h0975b: out <= 12'hfff;
      20'h0975c: out <= 12'hbbb;
      20'h0975d: out <= 12'h666;
      20'h0975e: out <= 12'h666;
      20'h0975f: out <= 12'h666;
      20'h09760: out <= 12'h000;
      20'h09761: out <= 12'h666;
      20'h09762: out <= 12'hfff;
      20'h09763: out <= 12'h666;
      20'h09764: out <= 12'hbbb;
      20'h09765: out <= 12'hfff;
      20'h09766: out <= 12'h666;
      20'h09767: out <= 12'h666;
      20'h09768: out <= 12'h666;
      20'h09769: out <= 12'h666;
      20'h0976a: out <= 12'h666;
      20'h0976b: out <= 12'hfff;
      20'h0976c: out <= 12'hbbb;
      20'h0976d: out <= 12'h666;
      20'h0976e: out <= 12'hfff;
      20'h0976f: out <= 12'h666;
      20'h09770: out <= 12'h603;
      20'h09771: out <= 12'h603;
      20'h09772: out <= 12'h603;
      20'h09773: out <= 12'h603;
      20'h09774: out <= 12'hf87;
      20'h09775: out <= 12'hf87;
      20'h09776: out <= 12'h000;
      20'h09777: out <= 12'h000;
      20'h09778: out <= 12'hf87;
      20'h09779: out <= 12'hf87;
      20'h0977a: out <= 12'hf87;
      20'h0977b: out <= 12'h000;
      20'h0977c: out <= 12'h000;
      20'h0977d: out <= 12'h000;
      20'h0977e: out <= 12'h000;
      20'h0977f: out <= 12'hf87;
      20'h09780: out <= 12'hf87;
      20'h09781: out <= 12'h000;
      20'h09782: out <= 12'h000;
      20'h09783: out <= 12'h000;
      20'h09784: out <= 12'h000;
      20'h09785: out <= 12'h000;
      20'h09786: out <= 12'h000;
      20'h09787: out <= 12'h000;
      20'h09788: out <= 12'h000;
      20'h09789: out <= 12'hf87;
      20'h0978a: out <= 12'hf87;
      20'h0978b: out <= 12'h000;
      20'h0978c: out <= 12'h000;
      20'h0978d: out <= 12'h000;
      20'h0978e: out <= 12'h000;
      20'h0978f: out <= 12'h000;
      20'h09790: out <= 12'h000;
      20'h09791: out <= 12'hf87;
      20'h09792: out <= 12'hf87;
      20'h09793: out <= 12'h000;
      20'h09794: out <= 12'h000;
      20'h09795: out <= 12'hf87;
      20'h09796: out <= 12'hf87;
      20'h09797: out <= 12'h000;
      20'h09798: out <= 12'hf87;
      20'h09799: out <= 12'hf87;
      20'h0979a: out <= 12'h000;
      20'h0979b: out <= 12'h000;
      20'h0979c: out <= 12'hf87;
      20'h0979d: out <= 12'hf87;
      20'h0979e: out <= 12'hf87;
      20'h0979f: out <= 12'hf87;
      20'h097a0: out <= 12'hf87;
      20'h097a1: out <= 12'hf87;
      20'h097a2: out <= 12'h000;
      20'h097a3: out <= 12'h000;
      20'h097a4: out <= 12'hf87;
      20'h097a5: out <= 12'hf87;
      20'h097a6: out <= 12'h000;
      20'h097a7: out <= 12'h000;
      20'h097a8: out <= 12'h000;
      20'h097a9: out <= 12'h000;
      20'h097aa: out <= 12'h000;
      20'h097ab: out <= 12'h000;
      20'h097ac: out <= 12'h000;
      20'h097ad: out <= 12'h000;
      20'h097ae: out <= 12'h000;
      20'h097af: out <= 12'h000;
      20'h097b0: out <= 12'hf87;
      20'h097b1: out <= 12'hf87;
      20'h097b2: out <= 12'h000;
      20'h097b3: out <= 12'h000;
      20'h097b4: out <= 12'hf87;
      20'h097b5: out <= 12'hf87;
      20'h097b6: out <= 12'h000;
      20'h097b7: out <= 12'h000;
      20'h097b8: out <= 12'h000;
      20'h097b9: out <= 12'hf87;
      20'h097ba: out <= 12'hf87;
      20'h097bb: out <= 12'h000;
      20'h097bc: out <= 12'hf87;
      20'h097bd: out <= 12'hf87;
      20'h097be: out <= 12'h000;
      20'h097bf: out <= 12'h000;
      20'h097c0: out <= 12'h000;
      20'h097c1: out <= 12'hf87;
      20'h097c2: out <= 12'hf87;
      20'h097c3: out <= 12'h000;
      20'h097c4: out <= 12'h603;
      20'h097c5: out <= 12'h603;
      20'h097c6: out <= 12'h603;
      20'h097c7: out <= 12'h603;
      20'h097c8: out <= 12'hee9;
      20'h097c9: out <= 12'hf87;
      20'h097ca: out <= 12'hee9;
      20'h097cb: out <= 12'hee9;
      20'h097cc: out <= 12'hee9;
      20'h097cd: out <= 12'hb27;
      20'h097ce: out <= 12'hf87;
      20'h097cf: out <= 12'hb27;
      20'h097d0: out <= 12'h000;
      20'h097d1: out <= 12'h000;
      20'h097d2: out <= 12'h000;
      20'h097d3: out <= 12'h000;
      20'h097d4: out <= 12'h000;
      20'h097d5: out <= 12'h000;
      20'h097d6: out <= 12'h000;
      20'h097d7: out <= 12'h000;
      20'h097d8: out <= 12'h000;
      20'h097d9: out <= 12'h000;
      20'h097da: out <= 12'h000;
      20'h097db: out <= 12'h000;
      20'h097dc: out <= 12'h000;
      20'h097dd: out <= 12'h000;
      20'h097de: out <= 12'h000;
      20'h097df: out <= 12'h72f;
      20'h097e0: out <= 12'hfff;
      20'h097e1: out <= 12'h72f;
      20'h097e2: out <= 12'h000;
      20'h097e3: out <= 12'h000;
      20'h097e4: out <= 12'h000;
      20'h097e5: out <= 12'h000;
      20'h097e6: out <= 12'h000;
      20'h097e7: out <= 12'h000;
      20'h097e8: out <= 12'h000;
      20'h097e9: out <= 12'h000;
      20'h097ea: out <= 12'h000;
      20'h097eb: out <= 12'h000;
      20'h097ec: out <= 12'h000;
      20'h097ed: out <= 12'h000;
      20'h097ee: out <= 12'h000;
      20'h097ef: out <= 12'h000;
      20'h097f0: out <= 12'h000;
      20'h097f1: out <= 12'h000;
      20'h097f2: out <= 12'h000;
      20'h097f3: out <= 12'h000;
      20'h097f4: out <= 12'h000;
      20'h097f5: out <= 12'h000;
      20'h097f6: out <= 12'h000;
      20'h097f7: out <= 12'h000;
      20'h097f8: out <= 12'h000;
      20'h097f9: out <= 12'h000;
      20'h097fa: out <= 12'h000;
      20'h097fb: out <= 12'h000;
      20'h097fc: out <= 12'h000;
      20'h097fd: out <= 12'h000;
      20'h097fe: out <= 12'h000;
      20'h097ff: out <= 12'h000;
      20'h09800: out <= 12'h000;
      20'h09801: out <= 12'h000;
      20'h09802: out <= 12'h000;
      20'h09803: out <= 12'h000;
      20'h09804: out <= 12'h000;
      20'h09805: out <= 12'h000;
      20'h09806: out <= 12'h000;
      20'h09807: out <= 12'h000;
      20'h09808: out <= 12'h222;
      20'h09809: out <= 12'h666;
      20'h0980a: out <= 12'h666;
      20'h0980b: out <= 12'h666;
      20'h0980c: out <= 12'hbbb;
      20'h0980d: out <= 12'hbbb;
      20'h0980e: out <= 12'hbbb;
      20'h0980f: out <= 12'hbbb;
      20'h09810: out <= 12'hbbb;
      20'h09811: out <= 12'hbbb;
      20'h09812: out <= 12'hbbb;
      20'h09813: out <= 12'h666;
      20'h09814: out <= 12'h666;
      20'h09815: out <= 12'h666;
      20'h09816: out <= 12'h666;
      20'h09817: out <= 12'h222;
      20'h09818: out <= 12'h000;
      20'h09819: out <= 12'h666;
      20'h0981a: out <= 12'h666;
      20'h0981b: out <= 12'h666;
      20'h0981c: out <= 12'hbbb;
      20'h0981d: out <= 12'hbbb;
      20'h0981e: out <= 12'hbbb;
      20'h0981f: out <= 12'hbbb;
      20'h09820: out <= 12'hbbb;
      20'h09821: out <= 12'hbbb;
      20'h09822: out <= 12'hbbb;
      20'h09823: out <= 12'h666;
      20'h09824: out <= 12'h666;
      20'h09825: out <= 12'h666;
      20'h09826: out <= 12'h666;
      20'h09827: out <= 12'h000;
      20'h09828: out <= 12'h222;
      20'h09829: out <= 12'h666;
      20'h0982a: out <= 12'h666;
      20'h0982b: out <= 12'h666;
      20'h0982c: out <= 12'hbbb;
      20'h0982d: out <= 12'hfff;
      20'h0982e: out <= 12'h666;
      20'h0982f: out <= 12'hfff;
      20'h09830: out <= 12'hfff;
      20'h09831: out <= 12'hfff;
      20'h09832: out <= 12'h666;
      20'h09833: out <= 12'hfff;
      20'h09834: out <= 12'hbbb;
      20'h09835: out <= 12'h666;
      20'h09836: out <= 12'h666;
      20'h09837: out <= 12'h666;
      20'h09838: out <= 12'h000;
      20'h09839: out <= 12'h666;
      20'h0983a: out <= 12'hfff;
      20'h0983b: out <= 12'h666;
      20'h0983c: out <= 12'hbbb;
      20'h0983d: out <= 12'hfff;
      20'h0983e: out <= 12'h666;
      20'h0983f: out <= 12'hbbb;
      20'h09840: out <= 12'hfff;
      20'h09841: out <= 12'hfff;
      20'h09842: out <= 12'h666;
      20'h09843: out <= 12'hfff;
      20'h09844: out <= 12'hbbb;
      20'h09845: out <= 12'h666;
      20'h09846: out <= 12'hfff;
      20'h09847: out <= 12'h666;
      20'h09848: out <= 12'h222;
      20'h09849: out <= 12'h666;
      20'h0984a: out <= 12'h666;
      20'h0984b: out <= 12'h666;
      20'h0984c: out <= 12'h666;
      20'h0984d: out <= 12'hbbb;
      20'h0984e: out <= 12'hbbb;
      20'h0984f: out <= 12'hbbb;
      20'h09850: out <= 12'hbbb;
      20'h09851: out <= 12'hbbb;
      20'h09852: out <= 12'hbbb;
      20'h09853: out <= 12'hbbb;
      20'h09854: out <= 12'h666;
      20'h09855: out <= 12'h666;
      20'h09856: out <= 12'h666;
      20'h09857: out <= 12'h222;
      20'h09858: out <= 12'h000;
      20'h09859: out <= 12'h666;
      20'h0985a: out <= 12'h666;
      20'h0985b: out <= 12'h666;
      20'h0985c: out <= 12'h666;
      20'h0985d: out <= 12'hbbb;
      20'h0985e: out <= 12'hbbb;
      20'h0985f: out <= 12'hbbb;
      20'h09860: out <= 12'hbbb;
      20'h09861: out <= 12'hbbb;
      20'h09862: out <= 12'hbbb;
      20'h09863: out <= 12'hbbb;
      20'h09864: out <= 12'h666;
      20'h09865: out <= 12'h666;
      20'h09866: out <= 12'h666;
      20'h09867: out <= 12'h000;
      20'h09868: out <= 12'h222;
      20'h09869: out <= 12'h666;
      20'h0986a: out <= 12'hfff;
      20'h0986b: out <= 12'h666;
      20'h0986c: out <= 12'h666;
      20'h0986d: out <= 12'hfff;
      20'h0986e: out <= 12'h666;
      20'h0986f: out <= 12'hbbb;
      20'h09870: out <= 12'hfff;
      20'h09871: out <= 12'hbbb;
      20'h09872: out <= 12'h666;
      20'h09873: out <= 12'hfff;
      20'h09874: out <= 12'h666;
      20'h09875: out <= 12'h666;
      20'h09876: out <= 12'hfff;
      20'h09877: out <= 12'h666;
      20'h09878: out <= 12'h000;
      20'h09879: out <= 12'h666;
      20'h0987a: out <= 12'h666;
      20'h0987b: out <= 12'h666;
      20'h0987c: out <= 12'h666;
      20'h0987d: out <= 12'hfff;
      20'h0987e: out <= 12'h666;
      20'h0987f: out <= 12'hbbb;
      20'h09880: out <= 12'hfff;
      20'h09881: out <= 12'hbbb;
      20'h09882: out <= 12'h666;
      20'h09883: out <= 12'hfff;
      20'h09884: out <= 12'h666;
      20'h09885: out <= 12'h666;
      20'h09886: out <= 12'h666;
      20'h09887: out <= 12'h666;
      20'h09888: out <= 12'h603;
      20'h09889: out <= 12'h603;
      20'h0988a: out <= 12'h603;
      20'h0988b: out <= 12'h603;
      20'h0988c: out <= 12'hf87;
      20'h0988d: out <= 12'hf87;
      20'h0988e: out <= 12'h000;
      20'h0988f: out <= 12'hf87;
      20'h09890: out <= 12'h000;
      20'h09891: out <= 12'hf87;
      20'h09892: out <= 12'hf87;
      20'h09893: out <= 12'h000;
      20'h09894: out <= 12'h000;
      20'h09895: out <= 12'h000;
      20'h09896: out <= 12'h000;
      20'h09897: out <= 12'hf87;
      20'h09898: out <= 12'hf87;
      20'h09899: out <= 12'h000;
      20'h0989a: out <= 12'h000;
      20'h0989b: out <= 12'h000;
      20'h0989c: out <= 12'h000;
      20'h0989d: out <= 12'h000;
      20'h0989e: out <= 12'h000;
      20'h0989f: out <= 12'hf87;
      20'h098a0: out <= 12'hf87;
      20'h098a1: out <= 12'hf87;
      20'h098a2: out <= 12'h000;
      20'h098a3: out <= 12'h000;
      20'h098a4: out <= 12'h000;
      20'h098a5: out <= 12'h000;
      20'h098a6: out <= 12'hf87;
      20'h098a7: out <= 12'hf87;
      20'h098a8: out <= 12'hf87;
      20'h098a9: out <= 12'hf87;
      20'h098aa: out <= 12'h000;
      20'h098ab: out <= 12'h000;
      20'h098ac: out <= 12'hf87;
      20'h098ad: out <= 12'hf87;
      20'h098ae: out <= 12'h000;
      20'h098af: out <= 12'h000;
      20'h098b0: out <= 12'hf87;
      20'h098b1: out <= 12'hf87;
      20'h098b2: out <= 12'h000;
      20'h098b3: out <= 12'h000;
      20'h098b4: out <= 12'h000;
      20'h098b5: out <= 12'h000;
      20'h098b6: out <= 12'h000;
      20'h098b7: out <= 12'h000;
      20'h098b8: out <= 12'h000;
      20'h098b9: out <= 12'hf87;
      20'h098ba: out <= 12'hf87;
      20'h098bb: out <= 12'h000;
      20'h098bc: out <= 12'hf87;
      20'h098bd: out <= 12'hf87;
      20'h098be: out <= 12'hf87;
      20'h098bf: out <= 12'hf87;
      20'h098c0: out <= 12'hf87;
      20'h098c1: out <= 12'hf87;
      20'h098c2: out <= 12'h000;
      20'h098c3: out <= 12'h000;
      20'h098c4: out <= 12'h000;
      20'h098c5: out <= 12'h000;
      20'h098c6: out <= 12'h000;
      20'h098c7: out <= 12'hf87;
      20'h098c8: out <= 12'hf87;
      20'h098c9: out <= 12'h000;
      20'h098ca: out <= 12'h000;
      20'h098cb: out <= 12'h000;
      20'h098cc: out <= 12'h000;
      20'h098cd: out <= 12'hf87;
      20'h098ce: out <= 12'hf87;
      20'h098cf: out <= 12'hf87;
      20'h098d0: out <= 12'hf87;
      20'h098d1: out <= 12'hf87;
      20'h098d2: out <= 12'h000;
      20'h098d3: out <= 12'h000;
      20'h098d4: out <= 12'h000;
      20'h098d5: out <= 12'hf87;
      20'h098d6: out <= 12'hf87;
      20'h098d7: out <= 12'hf87;
      20'h098d8: out <= 12'hf87;
      20'h098d9: out <= 12'hf87;
      20'h098da: out <= 12'hf87;
      20'h098db: out <= 12'h000;
      20'h098dc: out <= 12'h603;
      20'h098dd: out <= 12'h603;
      20'h098de: out <= 12'h603;
      20'h098df: out <= 12'h603;
      20'h098e0: out <= 12'hee9;
      20'h098e1: out <= 12'hf87;
      20'h098e2: out <= 12'hee9;
      20'h098e3: out <= 12'hf87;
      20'h098e4: out <= 12'hf87;
      20'h098e5: out <= 12'hb27;
      20'h098e6: out <= 12'hf87;
      20'h098e7: out <= 12'hb27;
      20'h098e8: out <= 12'h000;
      20'h098e9: out <= 12'h000;
      20'h098ea: out <= 12'h000;
      20'h098eb: out <= 12'h000;
      20'h098ec: out <= 12'h000;
      20'h098ed: out <= 12'h000;
      20'h098ee: out <= 12'h000;
      20'h098ef: out <= 12'h000;
      20'h098f0: out <= 12'h000;
      20'h098f1: out <= 12'hc7f;
      20'h098f2: out <= 12'h72f;
      20'h098f3: out <= 12'hc7f;
      20'h098f4: out <= 12'h000;
      20'h098f5: out <= 12'h000;
      20'h098f6: out <= 12'h000;
      20'h098f7: out <= 12'h72f;
      20'h098f8: out <= 12'hfff;
      20'h098f9: out <= 12'h72f;
      20'h098fa: out <= 12'h000;
      20'h098fb: out <= 12'h000;
      20'h098fc: out <= 12'h000;
      20'h098fd: out <= 12'hc7f;
      20'h098fe: out <= 12'h72f;
      20'h098ff: out <= 12'hc7f;
      20'h09900: out <= 12'h000;
      20'h09901: out <= 12'h000;
      20'h09902: out <= 12'h000;
      20'h09903: out <= 12'h000;
      20'h09904: out <= 12'h000;
      20'h09905: out <= 12'h000;
      20'h09906: out <= 12'h000;
      20'h09907: out <= 12'h000;
      20'h09908: out <= 12'h000;
      20'h09909: out <= 12'h000;
      20'h0990a: out <= 12'h000;
      20'h0990b: out <= 12'h000;
      20'h0990c: out <= 12'h000;
      20'h0990d: out <= 12'h000;
      20'h0990e: out <= 12'h000;
      20'h0990f: out <= 12'h000;
      20'h09910: out <= 12'h000;
      20'h09911: out <= 12'h000;
      20'h09912: out <= 12'h000;
      20'h09913: out <= 12'h000;
      20'h09914: out <= 12'h000;
      20'h09915: out <= 12'h000;
      20'h09916: out <= 12'h000;
      20'h09917: out <= 12'h000;
      20'h09918: out <= 12'h000;
      20'h09919: out <= 12'h000;
      20'h0991a: out <= 12'h000;
      20'h0991b: out <= 12'h000;
      20'h0991c: out <= 12'h000;
      20'h0991d: out <= 12'h000;
      20'h0991e: out <= 12'h000;
      20'h0991f: out <= 12'h000;
      20'h09920: out <= 12'h222;
      20'h09921: out <= 12'hbbb;
      20'h09922: out <= 12'hbbb;
      20'h09923: out <= 12'h666;
      20'h09924: out <= 12'h666;
      20'h09925: out <= 12'h666;
      20'h09926: out <= 12'h666;
      20'h09927: out <= 12'h666;
      20'h09928: out <= 12'h666;
      20'h09929: out <= 12'h666;
      20'h0992a: out <= 12'h666;
      20'h0992b: out <= 12'h666;
      20'h0992c: out <= 12'hbbb;
      20'h0992d: out <= 12'hbbb;
      20'h0992e: out <= 12'hbbb;
      20'h0992f: out <= 12'h222;
      20'h09930: out <= 12'h000;
      20'h09931: out <= 12'hbbb;
      20'h09932: out <= 12'hbbb;
      20'h09933: out <= 12'h666;
      20'h09934: out <= 12'h666;
      20'h09935: out <= 12'h666;
      20'h09936: out <= 12'h666;
      20'h09937: out <= 12'h666;
      20'h09938: out <= 12'h666;
      20'h09939: out <= 12'h666;
      20'h0993a: out <= 12'h666;
      20'h0993b: out <= 12'h666;
      20'h0993c: out <= 12'hbbb;
      20'h0993d: out <= 12'hbbb;
      20'h0993e: out <= 12'hbbb;
      20'h0993f: out <= 12'h000;
      20'h09940: out <= 12'h222;
      20'h09941: out <= 12'h666;
      20'h09942: out <= 12'hfff;
      20'h09943: out <= 12'h666;
      20'h09944: out <= 12'h666;
      20'h09945: out <= 12'hfff;
      20'h09946: out <= 12'h666;
      20'h09947: out <= 12'h666;
      20'h09948: out <= 12'h666;
      20'h09949: out <= 12'h666;
      20'h0994a: out <= 12'h666;
      20'h0994b: out <= 12'hfff;
      20'h0994c: out <= 12'h666;
      20'h0994d: out <= 12'h666;
      20'h0994e: out <= 12'hfff;
      20'h0994f: out <= 12'h666;
      20'h09950: out <= 12'h000;
      20'h09951: out <= 12'h666;
      20'h09952: out <= 12'h666;
      20'h09953: out <= 12'h666;
      20'h09954: out <= 12'h666;
      20'h09955: out <= 12'hfff;
      20'h09956: out <= 12'h666;
      20'h09957: out <= 12'h666;
      20'h09958: out <= 12'h666;
      20'h09959: out <= 12'h666;
      20'h0995a: out <= 12'h666;
      20'h0995b: out <= 12'hfff;
      20'h0995c: out <= 12'h666;
      20'h0995d: out <= 12'h666;
      20'h0995e: out <= 12'h666;
      20'h0995f: out <= 12'h666;
      20'h09960: out <= 12'h222;
      20'h09961: out <= 12'hbbb;
      20'h09962: out <= 12'hbbb;
      20'h09963: out <= 12'hbbb;
      20'h09964: out <= 12'h666;
      20'h09965: out <= 12'h666;
      20'h09966: out <= 12'h666;
      20'h09967: out <= 12'h666;
      20'h09968: out <= 12'h666;
      20'h09969: out <= 12'h666;
      20'h0996a: out <= 12'h666;
      20'h0996b: out <= 12'h666;
      20'h0996c: out <= 12'h666;
      20'h0996d: out <= 12'hbbb;
      20'h0996e: out <= 12'hbbb;
      20'h0996f: out <= 12'h222;
      20'h09970: out <= 12'h000;
      20'h09971: out <= 12'hbbb;
      20'h09972: out <= 12'hbbb;
      20'h09973: out <= 12'hbbb;
      20'h09974: out <= 12'h666;
      20'h09975: out <= 12'h666;
      20'h09976: out <= 12'h666;
      20'h09977: out <= 12'h666;
      20'h09978: out <= 12'h666;
      20'h09979: out <= 12'h666;
      20'h0997a: out <= 12'h666;
      20'h0997b: out <= 12'h666;
      20'h0997c: out <= 12'h666;
      20'h0997d: out <= 12'hbbb;
      20'h0997e: out <= 12'hbbb;
      20'h0997f: out <= 12'h000;
      20'h09980: out <= 12'h222;
      20'h09981: out <= 12'h666;
      20'h09982: out <= 12'h666;
      20'h09983: out <= 12'hbbb;
      20'h09984: out <= 12'h666;
      20'h09985: out <= 12'h666;
      20'h09986: out <= 12'h666;
      20'h09987: out <= 12'hbbb;
      20'h09988: out <= 12'hfff;
      20'h09989: out <= 12'hbbb;
      20'h0998a: out <= 12'h666;
      20'h0998b: out <= 12'h666;
      20'h0998c: out <= 12'h666;
      20'h0998d: out <= 12'hbbb;
      20'h0998e: out <= 12'h666;
      20'h0998f: out <= 12'h666;
      20'h09990: out <= 12'h000;
      20'h09991: out <= 12'h666;
      20'h09992: out <= 12'hfff;
      20'h09993: out <= 12'hbbb;
      20'h09994: out <= 12'h666;
      20'h09995: out <= 12'h666;
      20'h09996: out <= 12'h666;
      20'h09997: out <= 12'hbbb;
      20'h09998: out <= 12'hfff;
      20'h09999: out <= 12'hbbb;
      20'h0999a: out <= 12'h666;
      20'h0999b: out <= 12'h666;
      20'h0999c: out <= 12'h666;
      20'h0999d: out <= 12'hbbb;
      20'h0999e: out <= 12'hfff;
      20'h0999f: out <= 12'h666;
      20'h099a0: out <= 12'h603;
      20'h099a1: out <= 12'h603;
      20'h099a2: out <= 12'h603;
      20'h099a3: out <= 12'h603;
      20'h099a4: out <= 12'hf87;
      20'h099a5: out <= 12'hf87;
      20'h099a6: out <= 12'hf87;
      20'h099a7: out <= 12'h000;
      20'h099a8: out <= 12'h000;
      20'h099a9: out <= 12'hf87;
      20'h099aa: out <= 12'hf87;
      20'h099ab: out <= 12'h000;
      20'h099ac: out <= 12'h000;
      20'h099ad: out <= 12'h000;
      20'h099ae: out <= 12'h000;
      20'h099af: out <= 12'hf87;
      20'h099b0: out <= 12'hf87;
      20'h099b1: out <= 12'h000;
      20'h099b2: out <= 12'h000;
      20'h099b3: out <= 12'h000;
      20'h099b4: out <= 12'h000;
      20'h099b5: out <= 12'hf87;
      20'h099b6: out <= 12'hf87;
      20'h099b7: out <= 12'hf87;
      20'h099b8: out <= 12'h000;
      20'h099b9: out <= 12'h000;
      20'h099ba: out <= 12'h000;
      20'h099bb: out <= 12'h000;
      20'h099bc: out <= 12'h000;
      20'h099bd: out <= 12'h000;
      20'h099be: out <= 12'h000;
      20'h099bf: out <= 12'h000;
      20'h099c0: out <= 12'h000;
      20'h099c1: out <= 12'hf87;
      20'h099c2: out <= 12'hf87;
      20'h099c3: out <= 12'h000;
      20'h099c4: out <= 12'hf87;
      20'h099c5: out <= 12'hf87;
      20'h099c6: out <= 12'hf87;
      20'h099c7: out <= 12'hf87;
      20'h099c8: out <= 12'hf87;
      20'h099c9: out <= 12'hf87;
      20'h099ca: out <= 12'hf87;
      20'h099cb: out <= 12'h000;
      20'h099cc: out <= 12'h000;
      20'h099cd: out <= 12'h000;
      20'h099ce: out <= 12'h000;
      20'h099cf: out <= 12'h000;
      20'h099d0: out <= 12'h000;
      20'h099d1: out <= 12'hf87;
      20'h099d2: out <= 12'hf87;
      20'h099d3: out <= 12'h000;
      20'h099d4: out <= 12'hf87;
      20'h099d5: out <= 12'hf87;
      20'h099d6: out <= 12'h000;
      20'h099d7: out <= 12'h000;
      20'h099d8: out <= 12'h000;
      20'h099d9: out <= 12'hf87;
      20'h099da: out <= 12'hf87;
      20'h099db: out <= 12'h000;
      20'h099dc: out <= 12'h000;
      20'h099dd: out <= 12'h000;
      20'h099de: out <= 12'hf87;
      20'h099df: out <= 12'hf87;
      20'h099e0: out <= 12'h000;
      20'h099e1: out <= 12'h000;
      20'h099e2: out <= 12'h000;
      20'h099e3: out <= 12'h000;
      20'h099e4: out <= 12'hf87;
      20'h099e5: out <= 12'hf87;
      20'h099e6: out <= 12'h000;
      20'h099e7: out <= 12'h000;
      20'h099e8: out <= 12'h000;
      20'h099e9: out <= 12'hf87;
      20'h099ea: out <= 12'hf87;
      20'h099eb: out <= 12'h000;
      20'h099ec: out <= 12'h000;
      20'h099ed: out <= 12'h000;
      20'h099ee: out <= 12'h000;
      20'h099ef: out <= 12'h000;
      20'h099f0: out <= 12'h000;
      20'h099f1: out <= 12'hf87;
      20'h099f2: out <= 12'hf87;
      20'h099f3: out <= 12'h000;
      20'h099f4: out <= 12'h603;
      20'h099f5: out <= 12'h603;
      20'h099f6: out <= 12'h603;
      20'h099f7: out <= 12'h603;
      20'h099f8: out <= 12'hee9;
      20'h099f9: out <= 12'hf87;
      20'h099fa: out <= 12'hee9;
      20'h099fb: out <= 12'hf87;
      20'h099fc: out <= 12'hf87;
      20'h099fd: out <= 12'hb27;
      20'h099fe: out <= 12'hf87;
      20'h099ff: out <= 12'hb27;
      20'h09a00: out <= 12'h000;
      20'h09a01: out <= 12'h000;
      20'h09a02: out <= 12'h000;
      20'h09a03: out <= 12'h000;
      20'h09a04: out <= 12'h000;
      20'h09a05: out <= 12'h000;
      20'h09a06: out <= 12'h000;
      20'h09a07: out <= 12'h000;
      20'h09a08: out <= 12'h000;
      20'h09a09: out <= 12'hc7f;
      20'h09a0a: out <= 12'hfff;
      20'h09a0b: out <= 12'hc7f;
      20'h09a0c: out <= 12'h000;
      20'h09a0d: out <= 12'h72f;
      20'h09a0e: out <= 12'h72f;
      20'h09a0f: out <= 12'h72f;
      20'h09a10: out <= 12'hfff;
      20'h09a11: out <= 12'h72f;
      20'h09a12: out <= 12'h72f;
      20'h09a13: out <= 12'h72f;
      20'h09a14: out <= 12'h000;
      20'h09a15: out <= 12'hc7f;
      20'h09a16: out <= 12'hfff;
      20'h09a17: out <= 12'hc7f;
      20'h09a18: out <= 12'h000;
      20'h09a19: out <= 12'h000;
      20'h09a1a: out <= 12'h000;
      20'h09a1b: out <= 12'h000;
      20'h09a1c: out <= 12'h000;
      20'h09a1d: out <= 12'h000;
      20'h09a1e: out <= 12'h000;
      20'h09a1f: out <= 12'h000;
      20'h09a20: out <= 12'h000;
      20'h09a21: out <= 12'h000;
      20'h09a22: out <= 12'h000;
      20'h09a23: out <= 12'h000;
      20'h09a24: out <= 12'h000;
      20'h09a25: out <= 12'h000;
      20'h09a26: out <= 12'h000;
      20'h09a27: out <= 12'h000;
      20'h09a28: out <= 12'h000;
      20'h09a29: out <= 12'h000;
      20'h09a2a: out <= 12'h000;
      20'h09a2b: out <= 12'h000;
      20'h09a2c: out <= 12'h000;
      20'h09a2d: out <= 12'h000;
      20'h09a2e: out <= 12'h000;
      20'h09a2f: out <= 12'h000;
      20'h09a30: out <= 12'h000;
      20'h09a31: out <= 12'h000;
      20'h09a32: out <= 12'h000;
      20'h09a33: out <= 12'h000;
      20'h09a34: out <= 12'h000;
      20'h09a35: out <= 12'h000;
      20'h09a36: out <= 12'h000;
      20'h09a37: out <= 12'h000;
      20'h09a38: out <= 12'h222;
      20'h09a39: out <= 12'hfff;
      20'h09a3a: out <= 12'h666;
      20'h09a3b: out <= 12'hfff;
      20'h09a3c: out <= 12'h666;
      20'h09a3d: out <= 12'hfff;
      20'h09a3e: out <= 12'h666;
      20'h09a3f: out <= 12'hfff;
      20'h09a40: out <= 12'h666;
      20'h09a41: out <= 12'hfff;
      20'h09a42: out <= 12'h666;
      20'h09a43: out <= 12'hfff;
      20'h09a44: out <= 12'h666;
      20'h09a45: out <= 12'hfff;
      20'h09a46: out <= 12'h666;
      20'h09a47: out <= 12'h222;
      20'h09a48: out <= 12'h000;
      20'h09a49: out <= 12'h666;
      20'h09a4a: out <= 12'hfff;
      20'h09a4b: out <= 12'h666;
      20'h09a4c: out <= 12'hfff;
      20'h09a4d: out <= 12'h666;
      20'h09a4e: out <= 12'hfff;
      20'h09a4f: out <= 12'h666;
      20'h09a50: out <= 12'hfff;
      20'h09a51: out <= 12'h666;
      20'h09a52: out <= 12'hfff;
      20'h09a53: out <= 12'h666;
      20'h09a54: out <= 12'hfff;
      20'h09a55: out <= 12'h666;
      20'h09a56: out <= 12'hfff;
      20'h09a57: out <= 12'h000;
      20'h09a58: out <= 12'h222;
      20'h09a59: out <= 12'h666;
      20'h09a5a: out <= 12'h666;
      20'h09a5b: out <= 12'hbbb;
      20'h09a5c: out <= 12'h666;
      20'h09a5d: out <= 12'h666;
      20'h09a5e: out <= 12'hfff;
      20'h09a5f: out <= 12'hbbb;
      20'h09a60: out <= 12'h666;
      20'h09a61: out <= 12'hbbb;
      20'h09a62: out <= 12'hfff;
      20'h09a63: out <= 12'h666;
      20'h09a64: out <= 12'h666;
      20'h09a65: out <= 12'hbbb;
      20'h09a66: out <= 12'h666;
      20'h09a67: out <= 12'h666;
      20'h09a68: out <= 12'h000;
      20'h09a69: out <= 12'h666;
      20'h09a6a: out <= 12'hfff;
      20'h09a6b: out <= 12'hbbb;
      20'h09a6c: out <= 12'h666;
      20'h09a6d: out <= 12'h666;
      20'h09a6e: out <= 12'hfff;
      20'h09a6f: out <= 12'hbbb;
      20'h09a70: out <= 12'h666;
      20'h09a71: out <= 12'hbbb;
      20'h09a72: out <= 12'hfff;
      20'h09a73: out <= 12'h666;
      20'h09a74: out <= 12'h666;
      20'h09a75: out <= 12'hbbb;
      20'h09a76: out <= 12'hfff;
      20'h09a77: out <= 12'h666;
      20'h09a78: out <= 12'h222;
      20'h09a79: out <= 12'h666;
      20'h09a7a: out <= 12'hfff;
      20'h09a7b: out <= 12'h666;
      20'h09a7c: out <= 12'hfff;
      20'h09a7d: out <= 12'h666;
      20'h09a7e: out <= 12'hfff;
      20'h09a7f: out <= 12'h666;
      20'h09a80: out <= 12'hfff;
      20'h09a81: out <= 12'h666;
      20'h09a82: out <= 12'hfff;
      20'h09a83: out <= 12'h666;
      20'h09a84: out <= 12'hfff;
      20'h09a85: out <= 12'h666;
      20'h09a86: out <= 12'hfff;
      20'h09a87: out <= 12'h222;
      20'h09a88: out <= 12'h000;
      20'h09a89: out <= 12'hfff;
      20'h09a8a: out <= 12'h666;
      20'h09a8b: out <= 12'hfff;
      20'h09a8c: out <= 12'h666;
      20'h09a8d: out <= 12'hfff;
      20'h09a8e: out <= 12'h666;
      20'h09a8f: out <= 12'hfff;
      20'h09a90: out <= 12'h666;
      20'h09a91: out <= 12'hfff;
      20'h09a92: out <= 12'h666;
      20'h09a93: out <= 12'hfff;
      20'h09a94: out <= 12'h666;
      20'h09a95: out <= 12'hfff;
      20'h09a96: out <= 12'h666;
      20'h09a97: out <= 12'h000;
      20'h09a98: out <= 12'h222;
      20'h09a99: out <= 12'h666;
      20'h09a9a: out <= 12'hfff;
      20'h09a9b: out <= 12'hbbb;
      20'h09a9c: out <= 12'h666;
      20'h09a9d: out <= 12'h222;
      20'h09a9e: out <= 12'h222;
      20'h09a9f: out <= 12'hbbb;
      20'h09aa0: out <= 12'hfff;
      20'h09aa1: out <= 12'hbbb;
      20'h09aa2: out <= 12'h222;
      20'h09aa3: out <= 12'h222;
      20'h09aa4: out <= 12'h666;
      20'h09aa5: out <= 12'hbbb;
      20'h09aa6: out <= 12'hfff;
      20'h09aa7: out <= 12'h666;
      20'h09aa8: out <= 12'h000;
      20'h09aa9: out <= 12'h666;
      20'h09aaa: out <= 12'h666;
      20'h09aab: out <= 12'hbbb;
      20'h09aac: out <= 12'h666;
      20'h09aad: out <= 12'h000;
      20'h09aae: out <= 12'h000;
      20'h09aaf: out <= 12'hbbb;
      20'h09ab0: out <= 12'hfff;
      20'h09ab1: out <= 12'hbbb;
      20'h09ab2: out <= 12'h000;
      20'h09ab3: out <= 12'h000;
      20'h09ab4: out <= 12'h666;
      20'h09ab5: out <= 12'hbbb;
      20'h09ab6: out <= 12'h666;
      20'h09ab7: out <= 12'h666;
      20'h09ab8: out <= 12'h603;
      20'h09ab9: out <= 12'h603;
      20'h09aba: out <= 12'h603;
      20'h09abb: out <= 12'h603;
      20'h09abc: out <= 12'hf87;
      20'h09abd: out <= 12'hf87;
      20'h09abe: out <= 12'h000;
      20'h09abf: out <= 12'h000;
      20'h09ac0: out <= 12'h000;
      20'h09ac1: out <= 12'hf87;
      20'h09ac2: out <= 12'hf87;
      20'h09ac3: out <= 12'h000;
      20'h09ac4: out <= 12'h000;
      20'h09ac5: out <= 12'h000;
      20'h09ac6: out <= 12'h000;
      20'h09ac7: out <= 12'hf87;
      20'h09ac8: out <= 12'hf87;
      20'h09ac9: out <= 12'h000;
      20'h09aca: out <= 12'h000;
      20'h09acb: out <= 12'h000;
      20'h09acc: out <= 12'hf87;
      20'h09acd: out <= 12'hf87;
      20'h09ace: out <= 12'h000;
      20'h09acf: out <= 12'h000;
      20'h09ad0: out <= 12'h000;
      20'h09ad1: out <= 12'h000;
      20'h09ad2: out <= 12'h000;
      20'h09ad3: out <= 12'h000;
      20'h09ad4: out <= 12'hf87;
      20'h09ad5: out <= 12'hf87;
      20'h09ad6: out <= 12'h000;
      20'h09ad7: out <= 12'h000;
      20'h09ad8: out <= 12'h000;
      20'h09ad9: out <= 12'hf87;
      20'h09ada: out <= 12'hf87;
      20'h09adb: out <= 12'h000;
      20'h09adc: out <= 12'h000;
      20'h09add: out <= 12'h000;
      20'h09ade: out <= 12'h000;
      20'h09adf: out <= 12'h000;
      20'h09ae0: out <= 12'hf87;
      20'h09ae1: out <= 12'hf87;
      20'h09ae2: out <= 12'h000;
      20'h09ae3: out <= 12'h000;
      20'h09ae4: out <= 12'hf87;
      20'h09ae5: out <= 12'hf87;
      20'h09ae6: out <= 12'h000;
      20'h09ae7: out <= 12'h000;
      20'h09ae8: out <= 12'h000;
      20'h09ae9: out <= 12'hf87;
      20'h09aea: out <= 12'hf87;
      20'h09aeb: out <= 12'h000;
      20'h09aec: out <= 12'hf87;
      20'h09aed: out <= 12'hf87;
      20'h09aee: out <= 12'h000;
      20'h09aef: out <= 12'h000;
      20'h09af0: out <= 12'h000;
      20'h09af1: out <= 12'hf87;
      20'h09af2: out <= 12'hf87;
      20'h09af3: out <= 12'h000;
      20'h09af4: out <= 12'h000;
      20'h09af5: out <= 12'h000;
      20'h09af6: out <= 12'hf87;
      20'h09af7: out <= 12'hf87;
      20'h09af8: out <= 12'h000;
      20'h09af9: out <= 12'h000;
      20'h09afa: out <= 12'h000;
      20'h09afb: out <= 12'h000;
      20'h09afc: out <= 12'hf87;
      20'h09afd: out <= 12'hf87;
      20'h09afe: out <= 12'h000;
      20'h09aff: out <= 12'h000;
      20'h09b00: out <= 12'h000;
      20'h09b01: out <= 12'hf87;
      20'h09b02: out <= 12'hf87;
      20'h09b03: out <= 12'h000;
      20'h09b04: out <= 12'h000;
      20'h09b05: out <= 12'h000;
      20'h09b06: out <= 12'h000;
      20'h09b07: out <= 12'h000;
      20'h09b08: out <= 12'hf87;
      20'h09b09: out <= 12'hf87;
      20'h09b0a: out <= 12'h000;
      20'h09b0b: out <= 12'h000;
      20'h09b0c: out <= 12'h603;
      20'h09b0d: out <= 12'h603;
      20'h09b0e: out <= 12'h603;
      20'h09b0f: out <= 12'h603;
      20'h09b10: out <= 12'hee9;
      20'h09b11: out <= 12'hf87;
      20'h09b12: out <= 12'hee9;
      20'h09b13: out <= 12'hb27;
      20'h09b14: out <= 12'hb27;
      20'h09b15: out <= 12'hb27;
      20'h09b16: out <= 12'hf87;
      20'h09b17: out <= 12'hb27;
      20'h09b18: out <= 12'h000;
      20'h09b19: out <= 12'h000;
      20'h09b1a: out <= 12'h000;
      20'h09b1b: out <= 12'h000;
      20'h09b1c: out <= 12'h000;
      20'h09b1d: out <= 12'h000;
      20'h09b1e: out <= 12'h000;
      20'h09b1f: out <= 12'h000;
      20'h09b20: out <= 12'h000;
      20'h09b21: out <= 12'hc7f;
      20'h09b22: out <= 12'h72f;
      20'h09b23: out <= 12'h72f;
      20'h09b24: out <= 12'h72f;
      20'h09b25: out <= 12'hfff;
      20'h09b26: out <= 12'hc7f;
      20'h09b27: out <= 12'h72f;
      20'h09b28: out <= 12'h72f;
      20'h09b29: out <= 12'h72f;
      20'h09b2a: out <= 12'hc7f;
      20'h09b2b: out <= 12'hfff;
      20'h09b2c: out <= 12'h72f;
      20'h09b2d: out <= 12'h72f;
      20'h09b2e: out <= 12'h72f;
      20'h09b2f: out <= 12'hc7f;
      20'h09b30: out <= 12'h000;
      20'h09b31: out <= 12'h000;
      20'h09b32: out <= 12'h000;
      20'h09b33: out <= 12'h000;
      20'h09b34: out <= 12'h000;
      20'h09b35: out <= 12'h000;
      20'h09b36: out <= 12'h000;
      20'h09b37: out <= 12'h000;
      20'h09b38: out <= 12'h000;
      20'h09b39: out <= 12'h000;
      20'h09b3a: out <= 12'h000;
      20'h09b3b: out <= 12'h000;
      20'h09b3c: out <= 12'h000;
      20'h09b3d: out <= 12'h000;
      20'h09b3e: out <= 12'h000;
      20'h09b3f: out <= 12'h000;
      20'h09b40: out <= 12'h000;
      20'h09b41: out <= 12'h000;
      20'h09b42: out <= 12'h000;
      20'h09b43: out <= 12'h000;
      20'h09b44: out <= 12'h000;
      20'h09b45: out <= 12'h000;
      20'h09b46: out <= 12'h000;
      20'h09b47: out <= 12'h000;
      20'h09b48: out <= 12'h000;
      20'h09b49: out <= 12'h000;
      20'h09b4a: out <= 12'h000;
      20'h09b4b: out <= 12'h000;
      20'h09b4c: out <= 12'h000;
      20'h09b4d: out <= 12'h000;
      20'h09b4e: out <= 12'h000;
      20'h09b4f: out <= 12'h000;
      20'h09b50: out <= 12'h222;
      20'h09b51: out <= 12'h666;
      20'h09b52: out <= 12'h666;
      20'h09b53: out <= 12'h666;
      20'h09b54: out <= 12'h666;
      20'h09b55: out <= 12'h666;
      20'h09b56: out <= 12'h666;
      20'h09b57: out <= 12'h666;
      20'h09b58: out <= 12'h666;
      20'h09b59: out <= 12'h666;
      20'h09b5a: out <= 12'h666;
      20'h09b5b: out <= 12'h666;
      20'h09b5c: out <= 12'h666;
      20'h09b5d: out <= 12'h666;
      20'h09b5e: out <= 12'h666;
      20'h09b5f: out <= 12'h222;
      20'h09b60: out <= 12'h000;
      20'h09b61: out <= 12'h666;
      20'h09b62: out <= 12'h666;
      20'h09b63: out <= 12'h666;
      20'h09b64: out <= 12'h666;
      20'h09b65: out <= 12'h666;
      20'h09b66: out <= 12'h666;
      20'h09b67: out <= 12'h666;
      20'h09b68: out <= 12'h666;
      20'h09b69: out <= 12'h666;
      20'h09b6a: out <= 12'h666;
      20'h09b6b: out <= 12'h666;
      20'h09b6c: out <= 12'h666;
      20'h09b6d: out <= 12'h666;
      20'h09b6e: out <= 12'h666;
      20'h09b6f: out <= 12'h000;
      20'h09b70: out <= 12'h222;
      20'h09b71: out <= 12'h666;
      20'h09b72: out <= 12'hfff;
      20'h09b73: out <= 12'hbbb;
      20'h09b74: out <= 12'h666;
      20'h09b75: out <= 12'h222;
      20'h09b76: out <= 12'h666;
      20'h09b77: out <= 12'h666;
      20'h09b78: out <= 12'h666;
      20'h09b79: out <= 12'h666;
      20'h09b7a: out <= 12'h666;
      20'h09b7b: out <= 12'h222;
      20'h09b7c: out <= 12'h666;
      20'h09b7d: out <= 12'hbbb;
      20'h09b7e: out <= 12'hfff;
      20'h09b7f: out <= 12'h666;
      20'h09b80: out <= 12'h000;
      20'h09b81: out <= 12'h666;
      20'h09b82: out <= 12'h666;
      20'h09b83: out <= 12'hbbb;
      20'h09b84: out <= 12'h666;
      20'h09b85: out <= 12'h000;
      20'h09b86: out <= 12'h666;
      20'h09b87: out <= 12'h666;
      20'h09b88: out <= 12'h666;
      20'h09b89: out <= 12'h666;
      20'h09b8a: out <= 12'h666;
      20'h09b8b: out <= 12'h000;
      20'h09b8c: out <= 12'h666;
      20'h09b8d: out <= 12'hbbb;
      20'h09b8e: out <= 12'h666;
      20'h09b8f: out <= 12'h666;
      20'h09b90: out <= 12'h222;
      20'h09b91: out <= 12'h666;
      20'h09b92: out <= 12'h666;
      20'h09b93: out <= 12'h666;
      20'h09b94: out <= 12'h666;
      20'h09b95: out <= 12'h666;
      20'h09b96: out <= 12'h666;
      20'h09b97: out <= 12'h666;
      20'h09b98: out <= 12'h666;
      20'h09b99: out <= 12'h666;
      20'h09b9a: out <= 12'h666;
      20'h09b9b: out <= 12'h666;
      20'h09b9c: out <= 12'h666;
      20'h09b9d: out <= 12'h666;
      20'h09b9e: out <= 12'h666;
      20'h09b9f: out <= 12'h222;
      20'h09ba0: out <= 12'h000;
      20'h09ba1: out <= 12'h666;
      20'h09ba2: out <= 12'h666;
      20'h09ba3: out <= 12'h666;
      20'h09ba4: out <= 12'h666;
      20'h09ba5: out <= 12'h666;
      20'h09ba6: out <= 12'h666;
      20'h09ba7: out <= 12'h666;
      20'h09ba8: out <= 12'h666;
      20'h09ba9: out <= 12'h666;
      20'h09baa: out <= 12'h666;
      20'h09bab: out <= 12'h666;
      20'h09bac: out <= 12'h666;
      20'h09bad: out <= 12'h666;
      20'h09bae: out <= 12'h666;
      20'h09baf: out <= 12'h000;
      20'h09bb0: out <= 12'h222;
      20'h09bb1: out <= 12'h666;
      20'h09bb2: out <= 12'h666;
      20'h09bb3: out <= 12'hbbb;
      20'h09bb4: out <= 12'h666;
      20'h09bb5: out <= 12'h222;
      20'h09bb6: out <= 12'h222;
      20'h09bb7: out <= 12'hbbb;
      20'h09bb8: out <= 12'hfff;
      20'h09bb9: out <= 12'hbbb;
      20'h09bba: out <= 12'h222;
      20'h09bbb: out <= 12'h222;
      20'h09bbc: out <= 12'h666;
      20'h09bbd: out <= 12'hbbb;
      20'h09bbe: out <= 12'h666;
      20'h09bbf: out <= 12'h666;
      20'h09bc0: out <= 12'h000;
      20'h09bc1: out <= 12'h666;
      20'h09bc2: out <= 12'hfff;
      20'h09bc3: out <= 12'hbbb;
      20'h09bc4: out <= 12'h666;
      20'h09bc5: out <= 12'h000;
      20'h09bc6: out <= 12'h000;
      20'h09bc7: out <= 12'hbbb;
      20'h09bc8: out <= 12'hfff;
      20'h09bc9: out <= 12'hbbb;
      20'h09bca: out <= 12'h000;
      20'h09bcb: out <= 12'h000;
      20'h09bcc: out <= 12'h666;
      20'h09bcd: out <= 12'hbbb;
      20'h09bce: out <= 12'hfff;
      20'h09bcf: out <= 12'h666;
      20'h09bd0: out <= 12'h603;
      20'h09bd1: out <= 12'h603;
      20'h09bd2: out <= 12'h603;
      20'h09bd3: out <= 12'h603;
      20'h09bd4: out <= 12'h000;
      20'h09bd5: out <= 12'hf87;
      20'h09bd6: out <= 12'hf87;
      20'h09bd7: out <= 12'hf87;
      20'h09bd8: out <= 12'hf87;
      20'h09bd9: out <= 12'hf87;
      20'h09bda: out <= 12'h000;
      20'h09bdb: out <= 12'h000;
      20'h09bdc: out <= 12'h000;
      20'h09bdd: out <= 12'h000;
      20'h09bde: out <= 12'h000;
      20'h09bdf: out <= 12'hf87;
      20'h09be0: out <= 12'hf87;
      20'h09be1: out <= 12'h000;
      20'h09be2: out <= 12'h000;
      20'h09be3: out <= 12'h000;
      20'h09be4: out <= 12'hf87;
      20'h09be5: out <= 12'hf87;
      20'h09be6: out <= 12'hf87;
      20'h09be7: out <= 12'hf87;
      20'h09be8: out <= 12'hf87;
      20'h09be9: out <= 12'hf87;
      20'h09bea: out <= 12'hf87;
      20'h09beb: out <= 12'h000;
      20'h09bec: out <= 12'h000;
      20'h09bed: out <= 12'hf87;
      20'h09bee: out <= 12'hf87;
      20'h09bef: out <= 12'hf87;
      20'h09bf0: out <= 12'hf87;
      20'h09bf1: out <= 12'hf87;
      20'h09bf2: out <= 12'h000;
      20'h09bf3: out <= 12'h000;
      20'h09bf4: out <= 12'h000;
      20'h09bf5: out <= 12'h000;
      20'h09bf6: out <= 12'h000;
      20'h09bf7: out <= 12'h000;
      20'h09bf8: out <= 12'hf87;
      20'h09bf9: out <= 12'hf87;
      20'h09bfa: out <= 12'h000;
      20'h09bfb: out <= 12'h000;
      20'h09bfc: out <= 12'h000;
      20'h09bfd: out <= 12'hf87;
      20'h09bfe: out <= 12'hf87;
      20'h09bff: out <= 12'hf87;
      20'h09c00: out <= 12'hf87;
      20'h09c01: out <= 12'hf87;
      20'h09c02: out <= 12'h000;
      20'h09c03: out <= 12'h000;
      20'h09c04: out <= 12'h000;
      20'h09c05: out <= 12'hf87;
      20'h09c06: out <= 12'hf87;
      20'h09c07: out <= 12'hf87;
      20'h09c08: out <= 12'hf87;
      20'h09c09: out <= 12'hf87;
      20'h09c0a: out <= 12'h000;
      20'h09c0b: out <= 12'h000;
      20'h09c0c: out <= 12'h000;
      20'h09c0d: out <= 12'h000;
      20'h09c0e: out <= 12'hf87;
      20'h09c0f: out <= 12'hf87;
      20'h09c10: out <= 12'h000;
      20'h09c11: out <= 12'h000;
      20'h09c12: out <= 12'h000;
      20'h09c13: out <= 12'h000;
      20'h09c14: out <= 12'h000;
      20'h09c15: out <= 12'hf87;
      20'h09c16: out <= 12'hf87;
      20'h09c17: out <= 12'hf87;
      20'h09c18: out <= 12'hf87;
      20'h09c19: out <= 12'hf87;
      20'h09c1a: out <= 12'h000;
      20'h09c1b: out <= 12'h000;
      20'h09c1c: out <= 12'h000;
      20'h09c1d: out <= 12'hf87;
      20'h09c1e: out <= 12'hf87;
      20'h09c1f: out <= 12'hf87;
      20'h09c20: out <= 12'hf87;
      20'h09c21: out <= 12'h000;
      20'h09c22: out <= 12'h000;
      20'h09c23: out <= 12'h000;
      20'h09c24: out <= 12'h603;
      20'h09c25: out <= 12'h603;
      20'h09c26: out <= 12'h603;
      20'h09c27: out <= 12'h603;
      20'h09c28: out <= 12'hee9;
      20'h09c29: out <= 12'hf87;
      20'h09c2a: out <= 12'hf87;
      20'h09c2b: out <= 12'hf87;
      20'h09c2c: out <= 12'hf87;
      20'h09c2d: out <= 12'hf87;
      20'h09c2e: out <= 12'hf87;
      20'h09c2f: out <= 12'hb27;
      20'h09c30: out <= 12'h000;
      20'h09c31: out <= 12'h000;
      20'h09c32: out <= 12'h000;
      20'h09c33: out <= 12'h000;
      20'h09c34: out <= 12'h000;
      20'h09c35: out <= 12'h000;
      20'h09c36: out <= 12'h000;
      20'h09c37: out <= 12'h000;
      20'h09c38: out <= 12'h000;
      20'h09c39: out <= 12'hc7f;
      20'h09c3a: out <= 12'hfff;
      20'h09c3b: out <= 12'h72f;
      20'h09c3c: out <= 12'hfff;
      20'h09c3d: out <= 12'hc7f;
      20'h09c3e: out <= 12'h72f;
      20'h09c3f: out <= 12'h72f;
      20'h09c40: out <= 12'hc7f;
      20'h09c41: out <= 12'h72f;
      20'h09c42: out <= 12'h72f;
      20'h09c43: out <= 12'hc7f;
      20'h09c44: out <= 12'hfff;
      20'h09c45: out <= 12'h72f;
      20'h09c46: out <= 12'hfff;
      20'h09c47: out <= 12'hc7f;
      20'h09c48: out <= 12'h000;
      20'h09c49: out <= 12'h000;
      20'h09c4a: out <= 12'h000;
      20'h09c4b: out <= 12'h000;
      20'h09c4c: out <= 12'h000;
      20'h09c4d: out <= 12'h000;
      20'h09c4e: out <= 12'h000;
      20'h09c4f: out <= 12'h000;
      20'h09c50: out <= 12'h000;
      20'h09c51: out <= 12'h000;
      20'h09c52: out <= 12'h000;
      20'h09c53: out <= 12'h000;
      20'h09c54: out <= 12'h000;
      20'h09c55: out <= 12'h000;
      20'h09c56: out <= 12'h000;
      20'h09c57: out <= 12'h000;
      20'h09c58: out <= 12'h000;
      20'h09c59: out <= 12'h000;
      20'h09c5a: out <= 12'h000;
      20'h09c5b: out <= 12'h000;
      20'h09c5c: out <= 12'h000;
      20'h09c5d: out <= 12'h000;
      20'h09c5e: out <= 12'h000;
      20'h09c5f: out <= 12'h000;
      20'h09c60: out <= 12'h000;
      20'h09c61: out <= 12'h000;
      20'h09c62: out <= 12'h000;
      20'h09c63: out <= 12'h000;
      20'h09c64: out <= 12'h000;
      20'h09c65: out <= 12'h000;
      20'h09c66: out <= 12'h000;
      20'h09c67: out <= 12'h000;
      20'h09c68: out <= 12'h222;
      20'h09c69: out <= 12'h222;
      20'h09c6a: out <= 12'h222;
      20'h09c6b: out <= 12'h222;
      20'h09c6c: out <= 12'h222;
      20'h09c6d: out <= 12'h222;
      20'h09c6e: out <= 12'h222;
      20'h09c6f: out <= 12'h222;
      20'h09c70: out <= 12'h222;
      20'h09c71: out <= 12'h222;
      20'h09c72: out <= 12'h222;
      20'h09c73: out <= 12'h222;
      20'h09c74: out <= 12'h222;
      20'h09c75: out <= 12'h222;
      20'h09c76: out <= 12'h222;
      20'h09c77: out <= 12'h222;
      20'h09c78: out <= 12'h000;
      20'h09c79: out <= 12'h000;
      20'h09c7a: out <= 12'h000;
      20'h09c7b: out <= 12'h000;
      20'h09c7c: out <= 12'h000;
      20'h09c7d: out <= 12'h000;
      20'h09c7e: out <= 12'h000;
      20'h09c7f: out <= 12'h000;
      20'h09c80: out <= 12'h000;
      20'h09c81: out <= 12'h000;
      20'h09c82: out <= 12'h000;
      20'h09c83: out <= 12'h000;
      20'h09c84: out <= 12'h000;
      20'h09c85: out <= 12'h000;
      20'h09c86: out <= 12'h000;
      20'h09c87: out <= 12'h000;
      20'h09c88: out <= 12'h222;
      20'h09c89: out <= 12'h222;
      20'h09c8a: out <= 12'h222;
      20'h09c8b: out <= 12'h222;
      20'h09c8c: out <= 12'h222;
      20'h09c8d: out <= 12'h222;
      20'h09c8e: out <= 12'h222;
      20'h09c8f: out <= 12'h222;
      20'h09c90: out <= 12'h222;
      20'h09c91: out <= 12'h222;
      20'h09c92: out <= 12'h222;
      20'h09c93: out <= 12'h222;
      20'h09c94: out <= 12'h222;
      20'h09c95: out <= 12'h222;
      20'h09c96: out <= 12'h222;
      20'h09c97: out <= 12'h222;
      20'h09c98: out <= 12'h000;
      20'h09c99: out <= 12'h000;
      20'h09c9a: out <= 12'h000;
      20'h09c9b: out <= 12'h000;
      20'h09c9c: out <= 12'h000;
      20'h09c9d: out <= 12'h000;
      20'h09c9e: out <= 12'h000;
      20'h09c9f: out <= 12'h000;
      20'h09ca0: out <= 12'h000;
      20'h09ca1: out <= 12'h000;
      20'h09ca2: out <= 12'h000;
      20'h09ca3: out <= 12'h000;
      20'h09ca4: out <= 12'h000;
      20'h09ca5: out <= 12'h000;
      20'h09ca6: out <= 12'h000;
      20'h09ca7: out <= 12'h000;
      20'h09ca8: out <= 12'h222;
      20'h09ca9: out <= 12'h222;
      20'h09caa: out <= 12'h222;
      20'h09cab: out <= 12'h222;
      20'h09cac: out <= 12'h222;
      20'h09cad: out <= 12'h222;
      20'h09cae: out <= 12'h222;
      20'h09caf: out <= 12'h222;
      20'h09cb0: out <= 12'h222;
      20'h09cb1: out <= 12'h222;
      20'h09cb2: out <= 12'h222;
      20'h09cb3: out <= 12'h222;
      20'h09cb4: out <= 12'h222;
      20'h09cb5: out <= 12'h222;
      20'h09cb6: out <= 12'h222;
      20'h09cb7: out <= 12'h222;
      20'h09cb8: out <= 12'h000;
      20'h09cb9: out <= 12'h000;
      20'h09cba: out <= 12'h000;
      20'h09cbb: out <= 12'h000;
      20'h09cbc: out <= 12'h000;
      20'h09cbd: out <= 12'h000;
      20'h09cbe: out <= 12'h000;
      20'h09cbf: out <= 12'h000;
      20'h09cc0: out <= 12'h000;
      20'h09cc1: out <= 12'h000;
      20'h09cc2: out <= 12'h000;
      20'h09cc3: out <= 12'h000;
      20'h09cc4: out <= 12'h000;
      20'h09cc5: out <= 12'h000;
      20'h09cc6: out <= 12'h000;
      20'h09cc7: out <= 12'h000;
      20'h09cc8: out <= 12'h222;
      20'h09cc9: out <= 12'h222;
      20'h09cca: out <= 12'h222;
      20'h09ccb: out <= 12'h222;
      20'h09ccc: out <= 12'h222;
      20'h09ccd: out <= 12'h222;
      20'h09cce: out <= 12'hbbb;
      20'h09ccf: out <= 12'hbbb;
      20'h09cd0: out <= 12'hfff;
      20'h09cd1: out <= 12'hbbb;
      20'h09cd2: out <= 12'hbbb;
      20'h09cd3: out <= 12'h222;
      20'h09cd4: out <= 12'h222;
      20'h09cd5: out <= 12'h222;
      20'h09cd6: out <= 12'h222;
      20'h09cd7: out <= 12'h222;
      20'h09cd8: out <= 12'h000;
      20'h09cd9: out <= 12'h000;
      20'h09cda: out <= 12'h000;
      20'h09cdb: out <= 12'h000;
      20'h09cdc: out <= 12'h000;
      20'h09cdd: out <= 12'h000;
      20'h09cde: out <= 12'hbbb;
      20'h09cdf: out <= 12'hbbb;
      20'h09ce0: out <= 12'hfff;
      20'h09ce1: out <= 12'hbbb;
      20'h09ce2: out <= 12'hbbb;
      20'h09ce3: out <= 12'h000;
      20'h09ce4: out <= 12'h000;
      20'h09ce5: out <= 12'h000;
      20'h09ce6: out <= 12'h000;
      20'h09ce7: out <= 12'h000;
      20'h09ce8: out <= 12'h603;
      20'h09ce9: out <= 12'h603;
      20'h09cea: out <= 12'h603;
      20'h09ceb: out <= 12'h603;
      20'h09cec: out <= 12'h000;
      20'h09ced: out <= 12'h000;
      20'h09cee: out <= 12'h000;
      20'h09cef: out <= 12'h000;
      20'h09cf0: out <= 12'h000;
      20'h09cf1: out <= 12'h000;
      20'h09cf2: out <= 12'h000;
      20'h09cf3: out <= 12'h000;
      20'h09cf4: out <= 12'h000;
      20'h09cf5: out <= 12'h000;
      20'h09cf6: out <= 12'h000;
      20'h09cf7: out <= 12'h000;
      20'h09cf8: out <= 12'h000;
      20'h09cf9: out <= 12'h000;
      20'h09cfa: out <= 12'h000;
      20'h09cfb: out <= 12'h000;
      20'h09cfc: out <= 12'h000;
      20'h09cfd: out <= 12'h000;
      20'h09cfe: out <= 12'h000;
      20'h09cff: out <= 12'h000;
      20'h09d00: out <= 12'h000;
      20'h09d01: out <= 12'h000;
      20'h09d02: out <= 12'h000;
      20'h09d03: out <= 12'h000;
      20'h09d04: out <= 12'h000;
      20'h09d05: out <= 12'h000;
      20'h09d06: out <= 12'h000;
      20'h09d07: out <= 12'h000;
      20'h09d08: out <= 12'h000;
      20'h09d09: out <= 12'h000;
      20'h09d0a: out <= 12'h000;
      20'h09d0b: out <= 12'h000;
      20'h09d0c: out <= 12'h000;
      20'h09d0d: out <= 12'h000;
      20'h09d0e: out <= 12'h000;
      20'h09d0f: out <= 12'h000;
      20'h09d10: out <= 12'h000;
      20'h09d11: out <= 12'h000;
      20'h09d12: out <= 12'h000;
      20'h09d13: out <= 12'h000;
      20'h09d14: out <= 12'h000;
      20'h09d15: out <= 12'h000;
      20'h09d16: out <= 12'h000;
      20'h09d17: out <= 12'h000;
      20'h09d18: out <= 12'h000;
      20'h09d19: out <= 12'h000;
      20'h09d1a: out <= 12'h000;
      20'h09d1b: out <= 12'h000;
      20'h09d1c: out <= 12'h000;
      20'h09d1d: out <= 12'h000;
      20'h09d1e: out <= 12'h000;
      20'h09d1f: out <= 12'h000;
      20'h09d20: out <= 12'h000;
      20'h09d21: out <= 12'h000;
      20'h09d22: out <= 12'h000;
      20'h09d23: out <= 12'h000;
      20'h09d24: out <= 12'h000;
      20'h09d25: out <= 12'h000;
      20'h09d26: out <= 12'h000;
      20'h09d27: out <= 12'h000;
      20'h09d28: out <= 12'h000;
      20'h09d29: out <= 12'h000;
      20'h09d2a: out <= 12'h000;
      20'h09d2b: out <= 12'h000;
      20'h09d2c: out <= 12'h000;
      20'h09d2d: out <= 12'h000;
      20'h09d2e: out <= 12'h000;
      20'h09d2f: out <= 12'h000;
      20'h09d30: out <= 12'h000;
      20'h09d31: out <= 12'h000;
      20'h09d32: out <= 12'h000;
      20'h09d33: out <= 12'h000;
      20'h09d34: out <= 12'h000;
      20'h09d35: out <= 12'h000;
      20'h09d36: out <= 12'h000;
      20'h09d37: out <= 12'h000;
      20'h09d38: out <= 12'h000;
      20'h09d39: out <= 12'h000;
      20'h09d3a: out <= 12'h000;
      20'h09d3b: out <= 12'h000;
      20'h09d3c: out <= 12'h603;
      20'h09d3d: out <= 12'h603;
      20'h09d3e: out <= 12'h603;
      20'h09d3f: out <= 12'h603;
      20'h09d40: out <= 12'hb27;
      20'h09d41: out <= 12'hb27;
      20'h09d42: out <= 12'hb27;
      20'h09d43: out <= 12'hb27;
      20'h09d44: out <= 12'hb27;
      20'h09d45: out <= 12'hb27;
      20'h09d46: out <= 12'hb27;
      20'h09d47: out <= 12'hb27;
      20'h09d48: out <= 12'h000;
      20'h09d49: out <= 12'h000;
      20'h09d4a: out <= 12'h000;
      20'h09d4b: out <= 12'h000;
      20'h09d4c: out <= 12'h000;
      20'h09d4d: out <= 12'h000;
      20'h09d4e: out <= 12'h000;
      20'h09d4f: out <= 12'h000;
      20'h09d50: out <= 12'h000;
      20'h09d51: out <= 12'hc7f;
      20'h09d52: out <= 12'h72f;
      20'h09d53: out <= 12'h72f;
      20'h09d54: out <= 12'hc7f;
      20'h09d55: out <= 12'h72f;
      20'h09d56: out <= 12'h72f;
      20'h09d57: out <= 12'hc7f;
      20'h09d58: out <= 12'hfff;
      20'h09d59: out <= 12'hc7f;
      20'h09d5a: out <= 12'h72f;
      20'h09d5b: out <= 12'h72f;
      20'h09d5c: out <= 12'hc7f;
      20'h09d5d: out <= 12'h72f;
      20'h09d5e: out <= 12'h72f;
      20'h09d5f: out <= 12'hc7f;
      20'h09d60: out <= 12'h000;
      20'h09d61: out <= 12'h000;
      20'h09d62: out <= 12'h000;
      20'h09d63: out <= 12'h000;
      20'h09d64: out <= 12'h000;
      20'h09d65: out <= 12'h000;
      20'h09d66: out <= 12'h000;
      20'h09d67: out <= 12'h000;
      20'h09d68: out <= 12'h000;
      20'h09d69: out <= 12'h000;
      20'h09d6a: out <= 12'h000;
      20'h09d6b: out <= 12'h000;
      20'h09d6c: out <= 12'h000;
      20'h09d6d: out <= 12'h000;
      20'h09d6e: out <= 12'h000;
      20'h09d6f: out <= 12'h000;
      20'h09d70: out <= 12'h000;
      20'h09d71: out <= 12'h000;
      20'h09d72: out <= 12'h000;
      20'h09d73: out <= 12'h000;
      20'h09d74: out <= 12'h000;
      20'h09d75: out <= 12'h000;
      20'h09d76: out <= 12'h000;
      20'h09d77: out <= 12'h000;
      20'h09d78: out <= 12'h000;
      20'h09d79: out <= 12'h000;
      20'h09d7a: out <= 12'h000;
      20'h09d7b: out <= 12'h000;
      20'h09d7c: out <= 12'h000;
      20'h09d7d: out <= 12'h000;
      20'h09d7e: out <= 12'h000;
      20'h09d7f: out <= 12'h000;
      20'h09d80: out <= 12'h000;
      20'h09d81: out <= 12'h660;
      20'h09d82: out <= 12'h660;
      20'h09d83: out <= 12'h660;
      20'h09d84: out <= 12'h660;
      20'h09d85: out <= 12'h660;
      20'h09d86: out <= 12'h660;
      20'h09d87: out <= 12'h660;
      20'h09d88: out <= 12'h660;
      20'h09d89: out <= 12'h660;
      20'h09d8a: out <= 12'h660;
      20'h09d8b: out <= 12'h660;
      20'h09d8c: out <= 12'h660;
      20'h09d8d: out <= 12'h660;
      20'h09d8e: out <= 12'h660;
      20'h09d8f: out <= 12'h000;
      20'h09d90: out <= 12'h222;
      20'h09d91: out <= 12'h660;
      20'h09d92: out <= 12'h660;
      20'h09d93: out <= 12'h660;
      20'h09d94: out <= 12'h660;
      20'h09d95: out <= 12'h660;
      20'h09d96: out <= 12'h660;
      20'h09d97: out <= 12'h660;
      20'h09d98: out <= 12'h660;
      20'h09d99: out <= 12'h660;
      20'h09d9a: out <= 12'h660;
      20'h09d9b: out <= 12'h660;
      20'h09d9c: out <= 12'h660;
      20'h09d9d: out <= 12'h660;
      20'h09d9e: out <= 12'h660;
      20'h09d9f: out <= 12'h222;
      20'h09da0: out <= 12'h000;
      20'h09da1: out <= 12'h000;
      20'h09da2: out <= 12'h000;
      20'h09da3: out <= 12'h000;
      20'h09da4: out <= 12'h000;
      20'h09da5: out <= 12'h000;
      20'h09da6: out <= 12'h000;
      20'h09da7: out <= 12'h660;
      20'h09da8: out <= 12'hee9;
      20'h09da9: out <= 12'hbb0;
      20'h09daa: out <= 12'h000;
      20'h09dab: out <= 12'h000;
      20'h09dac: out <= 12'h000;
      20'h09dad: out <= 12'h000;
      20'h09dae: out <= 12'h000;
      20'h09daf: out <= 12'h000;
      20'h09db0: out <= 12'h222;
      20'h09db1: out <= 12'h222;
      20'h09db2: out <= 12'h222;
      20'h09db3: out <= 12'h222;
      20'h09db4: out <= 12'h222;
      20'h09db5: out <= 12'h222;
      20'h09db6: out <= 12'h222;
      20'h09db7: out <= 12'h660;
      20'h09db8: out <= 12'hee9;
      20'h09db9: out <= 12'hbb0;
      20'h09dba: out <= 12'h222;
      20'h09dbb: out <= 12'h222;
      20'h09dbc: out <= 12'h222;
      20'h09dbd: out <= 12'h222;
      20'h09dbe: out <= 12'h222;
      20'h09dbf: out <= 12'h222;
      20'h09dc0: out <= 12'h000;
      20'h09dc1: out <= 12'h660;
      20'h09dc2: out <= 12'h660;
      20'h09dc3: out <= 12'h660;
      20'h09dc4: out <= 12'h660;
      20'h09dc5: out <= 12'h660;
      20'h09dc6: out <= 12'h660;
      20'h09dc7: out <= 12'h660;
      20'h09dc8: out <= 12'h660;
      20'h09dc9: out <= 12'h660;
      20'h09dca: out <= 12'h660;
      20'h09dcb: out <= 12'h660;
      20'h09dcc: out <= 12'h660;
      20'h09dcd: out <= 12'h660;
      20'h09dce: out <= 12'h660;
      20'h09dcf: out <= 12'h000;
      20'h09dd0: out <= 12'h222;
      20'h09dd1: out <= 12'h660;
      20'h09dd2: out <= 12'h660;
      20'h09dd3: out <= 12'h660;
      20'h09dd4: out <= 12'h660;
      20'h09dd5: out <= 12'h660;
      20'h09dd6: out <= 12'h660;
      20'h09dd7: out <= 12'h660;
      20'h09dd8: out <= 12'h660;
      20'h09dd9: out <= 12'h660;
      20'h09dda: out <= 12'h660;
      20'h09ddb: out <= 12'h660;
      20'h09ddc: out <= 12'h660;
      20'h09ddd: out <= 12'h660;
      20'h09dde: out <= 12'h660;
      20'h09ddf: out <= 12'h222;
      20'h09de0: out <= 12'h000;
      20'h09de1: out <= 12'h000;
      20'h09de2: out <= 12'h000;
      20'h09de3: out <= 12'h000;
      20'h09de4: out <= 12'h000;
      20'h09de5: out <= 12'h000;
      20'h09de6: out <= 12'h000;
      20'h09de7: out <= 12'h000;
      20'h09de8: out <= 12'h000;
      20'h09de9: out <= 12'h000;
      20'h09dea: out <= 12'h000;
      20'h09deb: out <= 12'h000;
      20'h09dec: out <= 12'h000;
      20'h09ded: out <= 12'h000;
      20'h09dee: out <= 12'h000;
      20'h09def: out <= 12'h000;
      20'h09df0: out <= 12'h222;
      20'h09df1: out <= 12'h222;
      20'h09df2: out <= 12'h222;
      20'h09df3: out <= 12'h222;
      20'h09df4: out <= 12'h222;
      20'h09df5: out <= 12'h222;
      20'h09df6: out <= 12'h222;
      20'h09df7: out <= 12'h222;
      20'h09df8: out <= 12'h222;
      20'h09df9: out <= 12'h222;
      20'h09dfa: out <= 12'h222;
      20'h09dfb: out <= 12'h222;
      20'h09dfc: out <= 12'h222;
      20'h09dfd: out <= 12'h222;
      20'h09dfe: out <= 12'h222;
      20'h09dff: out <= 12'h222;
      20'h09e00: out <= 12'h603;
      20'h09e01: out <= 12'h603;
      20'h09e02: out <= 12'h603;
      20'h09e03: out <= 12'h603;
      20'h09e04: out <= 12'h000;
      20'h09e05: out <= 12'h4cd;
      20'h09e06: out <= 12'h4cd;
      20'h09e07: out <= 12'h4cd;
      20'h09e08: out <= 12'h4cd;
      20'h09e09: out <= 12'h4cd;
      20'h09e0a: out <= 12'h000;
      20'h09e0b: out <= 12'h000;
      20'h09e0c: out <= 12'h000;
      20'h09e0d: out <= 12'h000;
      20'h09e0e: out <= 12'h000;
      20'h09e0f: out <= 12'h4cd;
      20'h09e10: out <= 12'h4cd;
      20'h09e11: out <= 12'h000;
      20'h09e12: out <= 12'h000;
      20'h09e13: out <= 12'h000;
      20'h09e14: out <= 12'h000;
      20'h09e15: out <= 12'h4cd;
      20'h09e16: out <= 12'h4cd;
      20'h09e17: out <= 12'h4cd;
      20'h09e18: out <= 12'h4cd;
      20'h09e19: out <= 12'h4cd;
      20'h09e1a: out <= 12'h000;
      20'h09e1b: out <= 12'h000;
      20'h09e1c: out <= 12'h000;
      20'h09e1d: out <= 12'h4cd;
      20'h09e1e: out <= 12'h4cd;
      20'h09e1f: out <= 12'h4cd;
      20'h09e20: out <= 12'h4cd;
      20'h09e21: out <= 12'h4cd;
      20'h09e22: out <= 12'h000;
      20'h09e23: out <= 12'h000;
      20'h09e24: out <= 12'h000;
      20'h09e25: out <= 12'h000;
      20'h09e26: out <= 12'h000;
      20'h09e27: out <= 12'h4cd;
      20'h09e28: out <= 12'h4cd;
      20'h09e29: out <= 12'h4cd;
      20'h09e2a: out <= 12'h000;
      20'h09e2b: out <= 12'h000;
      20'h09e2c: out <= 12'h4cd;
      20'h09e2d: out <= 12'h4cd;
      20'h09e2e: out <= 12'h4cd;
      20'h09e2f: out <= 12'h4cd;
      20'h09e30: out <= 12'h4cd;
      20'h09e31: out <= 12'h4cd;
      20'h09e32: out <= 12'h4cd;
      20'h09e33: out <= 12'h000;
      20'h09e34: out <= 12'h000;
      20'h09e35: out <= 12'h000;
      20'h09e36: out <= 12'h4cd;
      20'h09e37: out <= 12'h4cd;
      20'h09e38: out <= 12'h4cd;
      20'h09e39: out <= 12'h4cd;
      20'h09e3a: out <= 12'h000;
      20'h09e3b: out <= 12'h000;
      20'h09e3c: out <= 12'h4cd;
      20'h09e3d: out <= 12'h4cd;
      20'h09e3e: out <= 12'h4cd;
      20'h09e3f: out <= 12'h4cd;
      20'h09e40: out <= 12'h4cd;
      20'h09e41: out <= 12'h4cd;
      20'h09e42: out <= 12'h4cd;
      20'h09e43: out <= 12'h000;
      20'h09e44: out <= 12'h000;
      20'h09e45: out <= 12'h4cd;
      20'h09e46: out <= 12'h4cd;
      20'h09e47: out <= 12'h4cd;
      20'h09e48: out <= 12'h4cd;
      20'h09e49: out <= 12'h4cd;
      20'h09e4a: out <= 12'h000;
      20'h09e4b: out <= 12'h000;
      20'h09e4c: out <= 12'h000;
      20'h09e4d: out <= 12'h4cd;
      20'h09e4e: out <= 12'h4cd;
      20'h09e4f: out <= 12'h4cd;
      20'h09e50: out <= 12'h4cd;
      20'h09e51: out <= 12'h4cd;
      20'h09e52: out <= 12'h000;
      20'h09e53: out <= 12'h000;
      20'h09e54: out <= 12'h603;
      20'h09e55: out <= 12'h603;
      20'h09e56: out <= 12'h603;
      20'h09e57: out <= 12'h603;
      20'h09e58: out <= 12'hee9;
      20'h09e59: out <= 12'hee9;
      20'h09e5a: out <= 12'hee9;
      20'h09e5b: out <= 12'hee9;
      20'h09e5c: out <= 12'hee9;
      20'h09e5d: out <= 12'hee9;
      20'h09e5e: out <= 12'hee9;
      20'h09e5f: out <= 12'hb27;
      20'h09e60: out <= 12'h000;
      20'h09e61: out <= 12'h000;
      20'h09e62: out <= 12'h000;
      20'h09e63: out <= 12'h000;
      20'h09e64: out <= 12'h000;
      20'h09e65: out <= 12'h000;
      20'h09e66: out <= 12'h000;
      20'h09e67: out <= 12'h000;
      20'h09e68: out <= 12'h000;
      20'h09e69: out <= 12'hc7f;
      20'h09e6a: out <= 12'hfff;
      20'h09e6b: out <= 12'h72f;
      20'h09e6c: out <= 12'hc7f;
      20'h09e6d: out <= 12'h72f;
      20'h09e6e: out <= 12'hc7f;
      20'h09e6f: out <= 12'hfff;
      20'h09e70: out <= 12'hfff;
      20'h09e71: out <= 12'hfff;
      20'h09e72: out <= 12'hc7f;
      20'h09e73: out <= 12'h72f;
      20'h09e74: out <= 12'hc7f;
      20'h09e75: out <= 12'h72f;
      20'h09e76: out <= 12'hfff;
      20'h09e77: out <= 12'hc7f;
      20'h09e78: out <= 12'h000;
      20'h09e79: out <= 12'h000;
      20'h09e7a: out <= 12'h000;
      20'h09e7b: out <= 12'h000;
      20'h09e7c: out <= 12'h000;
      20'h09e7d: out <= 12'h000;
      20'h09e7e: out <= 12'h000;
      20'h09e7f: out <= 12'h000;
      20'h09e80: out <= 12'h4cd;
      20'h09e81: out <= 12'h4cd;
      20'h09e82: out <= 12'h4cd;
      20'h09e83: out <= 12'h4cd;
      20'h09e84: out <= 12'h4cd;
      20'h09e85: out <= 12'h4cd;
      20'h09e86: out <= 12'h4cd;
      20'h09e87: out <= 12'h4cd;
      20'h09e88: out <= 12'h5ef;
      20'h09e89: out <= 12'h5ef;
      20'h09e8a: out <= 12'h5ef;
      20'h09e8b: out <= 12'h5ef;
      20'h09e8c: out <= 12'h5ef;
      20'h09e8d: out <= 12'h5ef;
      20'h09e8e: out <= 12'h5ef;
      20'h09e8f: out <= 12'h5ef;
      20'h09e90: out <= 12'h000;
      20'h09e91: out <= 12'h000;
      20'h09e92: out <= 12'h000;
      20'h09e93: out <= 12'h000;
      20'h09e94: out <= 12'h000;
      20'h09e95: out <= 12'h000;
      20'h09e96: out <= 12'h000;
      20'h09e97: out <= 12'h000;
      20'h09e98: out <= 12'h000;
      20'h09e99: out <= 12'hee9;
      20'h09e9a: out <= 12'h660;
      20'h09e9b: out <= 12'hee9;
      20'h09e9c: out <= 12'h660;
      20'h09e9d: out <= 12'hee9;
      20'h09e9e: out <= 12'h660;
      20'h09e9f: out <= 12'hee9;
      20'h09ea0: out <= 12'h660;
      20'h09ea1: out <= 12'hee9;
      20'h09ea2: out <= 12'h660;
      20'h09ea3: out <= 12'hee9;
      20'h09ea4: out <= 12'h660;
      20'h09ea5: out <= 12'hee9;
      20'h09ea6: out <= 12'h660;
      20'h09ea7: out <= 12'h000;
      20'h09ea8: out <= 12'h222;
      20'h09ea9: out <= 12'h660;
      20'h09eaa: out <= 12'hee9;
      20'h09eab: out <= 12'h660;
      20'h09eac: out <= 12'hee9;
      20'h09ead: out <= 12'h660;
      20'h09eae: out <= 12'hee9;
      20'h09eaf: out <= 12'h660;
      20'h09eb0: out <= 12'hee9;
      20'h09eb1: out <= 12'h660;
      20'h09eb2: out <= 12'hee9;
      20'h09eb3: out <= 12'h660;
      20'h09eb4: out <= 12'hee9;
      20'h09eb5: out <= 12'h660;
      20'h09eb6: out <= 12'hee9;
      20'h09eb7: out <= 12'h222;
      20'h09eb8: out <= 12'h000;
      20'h09eb9: out <= 12'h660;
      20'h09eba: out <= 12'h660;
      20'h09ebb: out <= 12'hbb0;
      20'h09ebc: out <= 12'h000;
      20'h09ebd: out <= 12'hbb0;
      20'h09ebe: out <= 12'hee9;
      20'h09ebf: out <= 12'h660;
      20'h09ec0: out <= 12'hee9;
      20'h09ec1: out <= 12'hbb0;
      20'h09ec2: out <= 12'h660;
      20'h09ec3: out <= 12'h660;
      20'h09ec4: out <= 12'h000;
      20'h09ec5: out <= 12'hbb0;
      20'h09ec6: out <= 12'hee9;
      20'h09ec7: out <= 12'h660;
      20'h09ec8: out <= 12'h222;
      20'h09ec9: out <= 12'h660;
      20'h09eca: out <= 12'hee9;
      20'h09ecb: out <= 12'hbb0;
      20'h09ecc: out <= 12'h222;
      20'h09ecd: out <= 12'hbb0;
      20'h09ece: out <= 12'hee9;
      20'h09ecf: out <= 12'h660;
      20'h09ed0: out <= 12'hee9;
      20'h09ed1: out <= 12'hbb0;
      20'h09ed2: out <= 12'h660;
      20'h09ed3: out <= 12'h660;
      20'h09ed4: out <= 12'h222;
      20'h09ed5: out <= 12'hbb0;
      20'h09ed6: out <= 12'h660;
      20'h09ed7: out <= 12'h660;
      20'h09ed8: out <= 12'h000;
      20'h09ed9: out <= 12'h660;
      20'h09eda: out <= 12'hee9;
      20'h09edb: out <= 12'h660;
      20'h09edc: out <= 12'hee9;
      20'h09edd: out <= 12'h660;
      20'h09ede: out <= 12'hee9;
      20'h09edf: out <= 12'h660;
      20'h09ee0: out <= 12'hee9;
      20'h09ee1: out <= 12'h660;
      20'h09ee2: out <= 12'hee9;
      20'h09ee3: out <= 12'h660;
      20'h09ee4: out <= 12'hee9;
      20'h09ee5: out <= 12'h660;
      20'h09ee6: out <= 12'hee9;
      20'h09ee7: out <= 12'h000;
      20'h09ee8: out <= 12'h222;
      20'h09ee9: out <= 12'hee9;
      20'h09eea: out <= 12'h660;
      20'h09eeb: out <= 12'hee9;
      20'h09eec: out <= 12'h660;
      20'h09eed: out <= 12'hee9;
      20'h09eee: out <= 12'h660;
      20'h09eef: out <= 12'hee9;
      20'h09ef0: out <= 12'h660;
      20'h09ef1: out <= 12'hee9;
      20'h09ef2: out <= 12'h660;
      20'h09ef3: out <= 12'hee9;
      20'h09ef4: out <= 12'h660;
      20'h09ef5: out <= 12'hee9;
      20'h09ef6: out <= 12'h660;
      20'h09ef7: out <= 12'h222;
      20'h09ef8: out <= 12'h000;
      20'h09ef9: out <= 12'h660;
      20'h09efa: out <= 12'hee9;
      20'h09efb: out <= 12'hbb0;
      20'h09efc: out <= 12'h000;
      20'h09efd: out <= 12'hee9;
      20'h09efe: out <= 12'hee9;
      20'h09eff: out <= 12'h660;
      20'h09f00: out <= 12'h660;
      20'h09f01: out <= 12'h660;
      20'h09f02: out <= 12'h660;
      20'h09f03: out <= 12'h660;
      20'h09f04: out <= 12'h000;
      20'h09f05: out <= 12'hbb0;
      20'h09f06: out <= 12'h660;
      20'h09f07: out <= 12'h660;
      20'h09f08: out <= 12'h222;
      20'h09f09: out <= 12'h660;
      20'h09f0a: out <= 12'h660;
      20'h09f0b: out <= 12'hbb0;
      20'h09f0c: out <= 12'h222;
      20'h09f0d: out <= 12'hee9;
      20'h09f0e: out <= 12'hee9;
      20'h09f0f: out <= 12'h660;
      20'h09f10: out <= 12'h660;
      20'h09f11: out <= 12'h660;
      20'h09f12: out <= 12'h660;
      20'h09f13: out <= 12'h660;
      20'h09f14: out <= 12'h222;
      20'h09f15: out <= 12'hbb0;
      20'h09f16: out <= 12'hee9;
      20'h09f17: out <= 12'h660;
      20'h09f18: out <= 12'h603;
      20'h09f19: out <= 12'h603;
      20'h09f1a: out <= 12'h603;
      20'h09f1b: out <= 12'h603;
      20'h09f1c: out <= 12'h4cd;
      20'h09f1d: out <= 12'h4cd;
      20'h09f1e: out <= 12'h000;
      20'h09f1f: out <= 12'h000;
      20'h09f20: out <= 12'h000;
      20'h09f21: out <= 12'h4cd;
      20'h09f22: out <= 12'h4cd;
      20'h09f23: out <= 12'h000;
      20'h09f24: out <= 12'h000;
      20'h09f25: out <= 12'h000;
      20'h09f26: out <= 12'h4cd;
      20'h09f27: out <= 12'h4cd;
      20'h09f28: out <= 12'h4cd;
      20'h09f29: out <= 12'h000;
      20'h09f2a: out <= 12'h000;
      20'h09f2b: out <= 12'h000;
      20'h09f2c: out <= 12'h4cd;
      20'h09f2d: out <= 12'h4cd;
      20'h09f2e: out <= 12'h000;
      20'h09f2f: out <= 12'h000;
      20'h09f30: out <= 12'h000;
      20'h09f31: out <= 12'h4cd;
      20'h09f32: out <= 12'h4cd;
      20'h09f33: out <= 12'h000;
      20'h09f34: out <= 12'h4cd;
      20'h09f35: out <= 12'h4cd;
      20'h09f36: out <= 12'h000;
      20'h09f37: out <= 12'h000;
      20'h09f38: out <= 12'h000;
      20'h09f39: out <= 12'h4cd;
      20'h09f3a: out <= 12'h4cd;
      20'h09f3b: out <= 12'h000;
      20'h09f3c: out <= 12'h000;
      20'h09f3d: out <= 12'h000;
      20'h09f3e: out <= 12'h4cd;
      20'h09f3f: out <= 12'h4cd;
      20'h09f40: out <= 12'h4cd;
      20'h09f41: out <= 12'h4cd;
      20'h09f42: out <= 12'h000;
      20'h09f43: out <= 12'h000;
      20'h09f44: out <= 12'h4cd;
      20'h09f45: out <= 12'h4cd;
      20'h09f46: out <= 12'h000;
      20'h09f47: out <= 12'h000;
      20'h09f48: out <= 12'h000;
      20'h09f49: out <= 12'h000;
      20'h09f4a: out <= 12'h000;
      20'h09f4b: out <= 12'h000;
      20'h09f4c: out <= 12'h000;
      20'h09f4d: out <= 12'h4cd;
      20'h09f4e: out <= 12'h4cd;
      20'h09f4f: out <= 12'h000;
      20'h09f50: out <= 12'h000;
      20'h09f51: out <= 12'h000;
      20'h09f52: out <= 12'h000;
      20'h09f53: out <= 12'h000;
      20'h09f54: out <= 12'h4cd;
      20'h09f55: out <= 12'h4cd;
      20'h09f56: out <= 12'h000;
      20'h09f57: out <= 12'h000;
      20'h09f58: out <= 12'h000;
      20'h09f59: out <= 12'h4cd;
      20'h09f5a: out <= 12'h4cd;
      20'h09f5b: out <= 12'h000;
      20'h09f5c: out <= 12'h4cd;
      20'h09f5d: out <= 12'h4cd;
      20'h09f5e: out <= 12'h000;
      20'h09f5f: out <= 12'h000;
      20'h09f60: out <= 12'h000;
      20'h09f61: out <= 12'h4cd;
      20'h09f62: out <= 12'h4cd;
      20'h09f63: out <= 12'h000;
      20'h09f64: out <= 12'h4cd;
      20'h09f65: out <= 12'h4cd;
      20'h09f66: out <= 12'h000;
      20'h09f67: out <= 12'h000;
      20'h09f68: out <= 12'h000;
      20'h09f69: out <= 12'h4cd;
      20'h09f6a: out <= 12'h4cd;
      20'h09f6b: out <= 12'h000;
      20'h09f6c: out <= 12'h603;
      20'h09f6d: out <= 12'h603;
      20'h09f6e: out <= 12'h603;
      20'h09f6f: out <= 12'h603;
      20'h09f70: out <= 12'hee9;
      20'h09f71: out <= 12'hf87;
      20'h09f72: out <= 12'hf87;
      20'h09f73: out <= 12'hf87;
      20'h09f74: out <= 12'hf87;
      20'h09f75: out <= 12'hf87;
      20'h09f76: out <= 12'hf87;
      20'h09f77: out <= 12'hb27;
      20'h09f78: out <= 12'h000;
      20'h09f79: out <= 12'h000;
      20'h09f7a: out <= 12'h000;
      20'h09f7b: out <= 12'h000;
      20'h09f7c: out <= 12'h000;
      20'h09f7d: out <= 12'h000;
      20'h09f7e: out <= 12'h000;
      20'h09f7f: out <= 12'h000;
      20'h09f80: out <= 12'h000;
      20'h09f81: out <= 12'hc7f;
      20'h09f82: out <= 12'h72f;
      20'h09f83: out <= 12'h72f;
      20'h09f84: out <= 12'hc7f;
      20'h09f85: out <= 12'h72f;
      20'h09f86: out <= 12'h72f;
      20'h09f87: out <= 12'hc7f;
      20'h09f88: out <= 12'hfff;
      20'h09f89: out <= 12'hc7f;
      20'h09f8a: out <= 12'h72f;
      20'h09f8b: out <= 12'h72f;
      20'h09f8c: out <= 12'hc7f;
      20'h09f8d: out <= 12'h72f;
      20'h09f8e: out <= 12'h72f;
      20'h09f8f: out <= 12'hc7f;
      20'h09f90: out <= 12'h000;
      20'h09f91: out <= 12'h000;
      20'h09f92: out <= 12'h4cd;
      20'h09f93: out <= 12'h000;
      20'h09f94: out <= 12'h000;
      20'h09f95: out <= 12'h000;
      20'h09f96: out <= 12'h4cd;
      20'h09f97: out <= 12'h000;
      20'h09f98: out <= 12'h4cd;
      20'h09f99: out <= 12'h4cd;
      20'h09f9a: out <= 12'h4cd;
      20'h09f9b: out <= 12'h4cd;
      20'h09f9c: out <= 12'h4cd;
      20'h09f9d: out <= 12'h4cd;
      20'h09f9e: out <= 12'h4cd;
      20'h09f9f: out <= 12'h4cd;
      20'h09fa0: out <= 12'h5ef;
      20'h09fa1: out <= 12'h5ef;
      20'h09fa2: out <= 12'h5ef;
      20'h09fa3: out <= 12'h5ef;
      20'h09fa4: out <= 12'h5ef;
      20'h09fa5: out <= 12'h5ef;
      20'h09fa6: out <= 12'h5ef;
      20'h09fa7: out <= 12'h5ef;
      20'h09fa8: out <= 12'h000;
      20'h09fa9: out <= 12'h000;
      20'h09faa: out <= 12'h000;
      20'h09fab: out <= 12'h000;
      20'h09fac: out <= 12'h000;
      20'h09fad: out <= 12'h000;
      20'h09fae: out <= 12'h000;
      20'h09faf: out <= 12'h000;
      20'h09fb0: out <= 12'h088;
      20'h09fb1: out <= 12'h088;
      20'h09fb2: out <= 12'h088;
      20'h09fb3: out <= 12'h088;
      20'h09fb4: out <= 12'h088;
      20'h09fb5: out <= 12'h088;
      20'h09fb6: out <= 12'h088;
      20'h09fb7: out <= 12'h088;
      20'h09fb8: out <= 12'h088;
      20'h09fb9: out <= 12'h088;
      20'h09fba: out <= 12'h088;
      20'h09fbb: out <= 12'h088;
      20'h09fbc: out <= 12'h088;
      20'h09fbd: out <= 12'h088;
      20'h09fbe: out <= 12'h088;
      20'h09fbf: out <= 12'h088;
      20'h09fc0: out <= 12'h088;
      20'h09fc1: out <= 12'h088;
      20'h09fc2: out <= 12'h088;
      20'h09fc3: out <= 12'h088;
      20'h09fc4: out <= 12'h088;
      20'h09fc5: out <= 12'h088;
      20'h09fc6: out <= 12'h088;
      20'h09fc7: out <= 12'h088;
      20'h09fc8: out <= 12'h088;
      20'h09fc9: out <= 12'h088;
      20'h09fca: out <= 12'h088;
      20'h09fcb: out <= 12'h088;
      20'h09fcc: out <= 12'h088;
      20'h09fcd: out <= 12'h088;
      20'h09fce: out <= 12'h088;
      20'h09fcf: out <= 12'h088;
      20'h09fd0: out <= 12'h088;
      20'h09fd1: out <= 12'h088;
      20'h09fd2: out <= 12'h088;
      20'h09fd3: out <= 12'h088;
      20'h09fd4: out <= 12'h088;
      20'h09fd5: out <= 12'h088;
      20'h09fd6: out <= 12'h088;
      20'h09fd7: out <= 12'h088;
      20'h09fd8: out <= 12'h088;
      20'h09fd9: out <= 12'h088;
      20'h09fda: out <= 12'h088;
      20'h09fdb: out <= 12'h088;
      20'h09fdc: out <= 12'h088;
      20'h09fdd: out <= 12'h088;
      20'h09fde: out <= 12'h088;
      20'h09fdf: out <= 12'h088;
      20'h09fe0: out <= 12'h088;
      20'h09fe1: out <= 12'h088;
      20'h09fe2: out <= 12'h088;
      20'h09fe3: out <= 12'h088;
      20'h09fe4: out <= 12'h088;
      20'h09fe5: out <= 12'h088;
      20'h09fe6: out <= 12'h088;
      20'h09fe7: out <= 12'h088;
      20'h09fe8: out <= 12'h088;
      20'h09fe9: out <= 12'h088;
      20'h09fea: out <= 12'h088;
      20'h09feb: out <= 12'h088;
      20'h09fec: out <= 12'h088;
      20'h09fed: out <= 12'h088;
      20'h09fee: out <= 12'h088;
      20'h09fef: out <= 12'h088;
      20'h09ff0: out <= 12'h088;
      20'h09ff1: out <= 12'h088;
      20'h09ff2: out <= 12'h088;
      20'h09ff3: out <= 12'h088;
      20'h09ff4: out <= 12'h088;
      20'h09ff5: out <= 12'h088;
      20'h09ff6: out <= 12'h088;
      20'h09ff7: out <= 12'h088;
      20'h09ff8: out <= 12'h088;
      20'h09ff9: out <= 12'h088;
      20'h09ffa: out <= 12'h088;
      20'h09ffb: out <= 12'h088;
      20'h09ffc: out <= 12'h088;
      20'h09ffd: out <= 12'h088;
      20'h09ffe: out <= 12'h088;
      20'h09fff: out <= 12'h088;
      20'h0a000: out <= 12'h088;
      20'h0a001: out <= 12'h088;
      20'h0a002: out <= 12'h088;
      20'h0a003: out <= 12'h088;
      20'h0a004: out <= 12'h088;
      20'h0a005: out <= 12'h088;
      20'h0a006: out <= 12'h088;
      20'h0a007: out <= 12'h088;
      20'h0a008: out <= 12'h088;
      20'h0a009: out <= 12'h088;
      20'h0a00a: out <= 12'h088;
      20'h0a00b: out <= 12'h088;
      20'h0a00c: out <= 12'h088;
      20'h0a00d: out <= 12'h088;
      20'h0a00e: out <= 12'h088;
      20'h0a00f: out <= 12'h088;
      20'h0a010: out <= 12'h088;
      20'h0a011: out <= 12'h088;
      20'h0a012: out <= 12'h088;
      20'h0a013: out <= 12'h088;
      20'h0a014: out <= 12'h088;
      20'h0a015: out <= 12'h088;
      20'h0a016: out <= 12'h088;
      20'h0a017: out <= 12'h088;
      20'h0a018: out <= 12'h088;
      20'h0a019: out <= 12'hbb0;
      20'h0a01a: out <= 12'h660;
      20'h0a01b: out <= 12'h660;
      20'h0a01c: out <= 12'h660;
      20'h0a01d: out <= 12'hbb0;
      20'h0a01e: out <= 12'hee9;
      20'h0a01f: out <= 12'h660;
      20'h0a020: out <= 12'h222;
      20'h0a021: out <= 12'h660;
      20'h0a022: out <= 12'hee9;
      20'h0a023: out <= 12'hbb0;
      20'h0a024: out <= 12'hee9;
      20'h0a025: out <= 12'hee9;
      20'h0a026: out <= 12'hee9;
      20'h0a027: out <= 12'hbb0;
      20'h0a028: out <= 12'hbb0;
      20'h0a029: out <= 12'hbb0;
      20'h0a02a: out <= 12'h660;
      20'h0a02b: out <= 12'h660;
      20'h0a02c: out <= 12'h660;
      20'h0a02d: out <= 12'hbb0;
      20'h0a02e: out <= 12'h660;
      20'h0a02f: out <= 12'h660;
      20'h0a030: out <= 12'h603;
      20'h0a031: out <= 12'h603;
      20'h0a032: out <= 12'h603;
      20'h0a033: out <= 12'h603;
      20'h0a034: out <= 12'h4cd;
      20'h0a035: out <= 12'h4cd;
      20'h0a036: out <= 12'h000;
      20'h0a037: out <= 12'h000;
      20'h0a038: out <= 12'h4cd;
      20'h0a039: out <= 12'h4cd;
      20'h0a03a: out <= 12'h4cd;
      20'h0a03b: out <= 12'h000;
      20'h0a03c: out <= 12'h000;
      20'h0a03d: out <= 12'h000;
      20'h0a03e: out <= 12'h000;
      20'h0a03f: out <= 12'h4cd;
      20'h0a040: out <= 12'h4cd;
      20'h0a041: out <= 12'h000;
      20'h0a042: out <= 12'h000;
      20'h0a043: out <= 12'h000;
      20'h0a044: out <= 12'h000;
      20'h0a045: out <= 12'h000;
      20'h0a046: out <= 12'h000;
      20'h0a047: out <= 12'h000;
      20'h0a048: out <= 12'h000;
      20'h0a049: out <= 12'h4cd;
      20'h0a04a: out <= 12'h4cd;
      20'h0a04b: out <= 12'h000;
      20'h0a04c: out <= 12'h000;
      20'h0a04d: out <= 12'h000;
      20'h0a04e: out <= 12'h000;
      20'h0a04f: out <= 12'h000;
      20'h0a050: out <= 12'h000;
      20'h0a051: out <= 12'h4cd;
      20'h0a052: out <= 12'h4cd;
      20'h0a053: out <= 12'h000;
      20'h0a054: out <= 12'h000;
      20'h0a055: out <= 12'h4cd;
      20'h0a056: out <= 12'h4cd;
      20'h0a057: out <= 12'h000;
      20'h0a058: out <= 12'h4cd;
      20'h0a059: out <= 12'h4cd;
      20'h0a05a: out <= 12'h000;
      20'h0a05b: out <= 12'h000;
      20'h0a05c: out <= 12'h4cd;
      20'h0a05d: out <= 12'h4cd;
      20'h0a05e: out <= 12'h4cd;
      20'h0a05f: out <= 12'h4cd;
      20'h0a060: out <= 12'h4cd;
      20'h0a061: out <= 12'h4cd;
      20'h0a062: out <= 12'h000;
      20'h0a063: out <= 12'h000;
      20'h0a064: out <= 12'h4cd;
      20'h0a065: out <= 12'h4cd;
      20'h0a066: out <= 12'h000;
      20'h0a067: out <= 12'h000;
      20'h0a068: out <= 12'h000;
      20'h0a069: out <= 12'h000;
      20'h0a06a: out <= 12'h000;
      20'h0a06b: out <= 12'h000;
      20'h0a06c: out <= 12'h000;
      20'h0a06d: out <= 12'h000;
      20'h0a06e: out <= 12'h000;
      20'h0a06f: out <= 12'h000;
      20'h0a070: out <= 12'h4cd;
      20'h0a071: out <= 12'h4cd;
      20'h0a072: out <= 12'h000;
      20'h0a073: out <= 12'h000;
      20'h0a074: out <= 12'h4cd;
      20'h0a075: out <= 12'h4cd;
      20'h0a076: out <= 12'h000;
      20'h0a077: out <= 12'h000;
      20'h0a078: out <= 12'h000;
      20'h0a079: out <= 12'h4cd;
      20'h0a07a: out <= 12'h4cd;
      20'h0a07b: out <= 12'h000;
      20'h0a07c: out <= 12'h4cd;
      20'h0a07d: out <= 12'h4cd;
      20'h0a07e: out <= 12'h000;
      20'h0a07f: out <= 12'h000;
      20'h0a080: out <= 12'h000;
      20'h0a081: out <= 12'h4cd;
      20'h0a082: out <= 12'h4cd;
      20'h0a083: out <= 12'h000;
      20'h0a084: out <= 12'h603;
      20'h0a085: out <= 12'h603;
      20'h0a086: out <= 12'h603;
      20'h0a087: out <= 12'h603;
      20'h0a088: out <= 12'hee9;
      20'h0a089: out <= 12'hf87;
      20'h0a08a: out <= 12'hee9;
      20'h0a08b: out <= 12'hee9;
      20'h0a08c: out <= 12'hee9;
      20'h0a08d: out <= 12'hb27;
      20'h0a08e: out <= 12'hf87;
      20'h0a08f: out <= 12'hb27;
      20'h0a090: out <= 12'h000;
      20'h0a091: out <= 12'h000;
      20'h0a092: out <= 12'h000;
      20'h0a093: out <= 12'h000;
      20'h0a094: out <= 12'h000;
      20'h0a095: out <= 12'h000;
      20'h0a096: out <= 12'h000;
      20'h0a097: out <= 12'h000;
      20'h0a098: out <= 12'h000;
      20'h0a099: out <= 12'hc7f;
      20'h0a09a: out <= 12'hfff;
      20'h0a09b: out <= 12'h72f;
      20'h0a09c: out <= 12'hc7f;
      20'h0a09d: out <= 12'hc7f;
      20'h0a09e: out <= 12'h72f;
      20'h0a09f: out <= 12'h72f;
      20'h0a0a0: out <= 12'hc7f;
      20'h0a0a1: out <= 12'h72f;
      20'h0a0a2: out <= 12'h72f;
      20'h0a0a3: out <= 12'hc7f;
      20'h0a0a4: out <= 12'hc7f;
      20'h0a0a5: out <= 12'h72f;
      20'h0a0a6: out <= 12'hfff;
      20'h0a0a7: out <= 12'hc7f;
      20'h0a0a8: out <= 12'h000;
      20'h0a0a9: out <= 12'h000;
      20'h0a0aa: out <= 12'h000;
      20'h0a0ab: out <= 12'h4cd;
      20'h0a0ac: out <= 12'h000;
      20'h0a0ad: out <= 12'h4cd;
      20'h0a0ae: out <= 12'h000;
      20'h0a0af: out <= 12'h000;
      20'h0a0b0: out <= 12'h4cd;
      20'h0a0b1: out <= 12'h4cd;
      20'h0a0b2: out <= 12'h4cd;
      20'h0a0b3: out <= 12'h4cd;
      20'h0a0b4: out <= 12'h4cd;
      20'h0a0b5: out <= 12'h4cd;
      20'h0a0b6: out <= 12'h4cd;
      20'h0a0b7: out <= 12'h4cd;
      20'h0a0b8: out <= 12'h5ef;
      20'h0a0b9: out <= 12'h5ef;
      20'h0a0ba: out <= 12'h5ef;
      20'h0a0bb: out <= 12'h5ef;
      20'h0a0bc: out <= 12'h5ef;
      20'h0a0bd: out <= 12'h5ef;
      20'h0a0be: out <= 12'h5ef;
      20'h0a0bf: out <= 12'h5ef;
      20'h0a0c0: out <= 12'h000;
      20'h0a0c1: out <= 12'h000;
      20'h0a0c2: out <= 12'h000;
      20'h0a0c3: out <= 12'h000;
      20'h0a0c4: out <= 12'h000;
      20'h0a0c5: out <= 12'h000;
      20'h0a0c6: out <= 12'h000;
      20'h0a0c7: out <= 12'h000;
      20'h0a0c8: out <= 12'h088;
      20'h0a0c9: out <= 12'h088;
      20'h0a0ca: out <= 12'h088;
      20'h0a0cb: out <= 12'h088;
      20'h0a0cc: out <= 12'h088;
      20'h0a0cd: out <= 12'h088;
      20'h0a0ce: out <= 12'h088;
      20'h0a0cf: out <= 12'h088;
      20'h0a0d0: out <= 12'h088;
      20'h0a0d1: out <= 12'h088;
      20'h0a0d2: out <= 12'h088;
      20'h0a0d3: out <= 12'h088;
      20'h0a0d4: out <= 12'h088;
      20'h0a0d5: out <= 12'h088;
      20'h0a0d6: out <= 12'h088;
      20'h0a0d7: out <= 12'h088;
      20'h0a0d8: out <= 12'h088;
      20'h0a0d9: out <= 12'h088;
      20'h0a0da: out <= 12'h088;
      20'h0a0db: out <= 12'h088;
      20'h0a0dc: out <= 12'h088;
      20'h0a0dd: out <= 12'h088;
      20'h0a0de: out <= 12'h088;
      20'h0a0df: out <= 12'h088;
      20'h0a0e0: out <= 12'h088;
      20'h0a0e1: out <= 12'h088;
      20'h0a0e2: out <= 12'h088;
      20'h0a0e3: out <= 12'h088;
      20'h0a0e4: out <= 12'h088;
      20'h0a0e5: out <= 12'h088;
      20'h0a0e6: out <= 12'h088;
      20'h0a0e7: out <= 12'h088;
      20'h0a0e8: out <= 12'h088;
      20'h0a0e9: out <= 12'h088;
      20'h0a0ea: out <= 12'h088;
      20'h0a0eb: out <= 12'h088;
      20'h0a0ec: out <= 12'h088;
      20'h0a0ed: out <= 12'h088;
      20'h0a0ee: out <= 12'h088;
      20'h0a0ef: out <= 12'h088;
      20'h0a0f0: out <= 12'h088;
      20'h0a0f1: out <= 12'h088;
      20'h0a0f2: out <= 12'h088;
      20'h0a0f3: out <= 12'h088;
      20'h0a0f4: out <= 12'h088;
      20'h0a0f5: out <= 12'h088;
      20'h0a0f6: out <= 12'h088;
      20'h0a0f7: out <= 12'h088;
      20'h0a0f8: out <= 12'h088;
      20'h0a0f9: out <= 12'h088;
      20'h0a0fa: out <= 12'h088;
      20'h0a0fb: out <= 12'h088;
      20'h0a0fc: out <= 12'h088;
      20'h0a0fd: out <= 12'h088;
      20'h0a0fe: out <= 12'h088;
      20'h0a0ff: out <= 12'h088;
      20'h0a100: out <= 12'h088;
      20'h0a101: out <= 12'h088;
      20'h0a102: out <= 12'h088;
      20'h0a103: out <= 12'h088;
      20'h0a104: out <= 12'h088;
      20'h0a105: out <= 12'h088;
      20'h0a106: out <= 12'h088;
      20'h0a107: out <= 12'h088;
      20'h0a108: out <= 12'h088;
      20'h0a109: out <= 12'h088;
      20'h0a10a: out <= 12'h088;
      20'h0a10b: out <= 12'h088;
      20'h0a10c: out <= 12'h088;
      20'h0a10d: out <= 12'h088;
      20'h0a10e: out <= 12'h088;
      20'h0a10f: out <= 12'h088;
      20'h0a110: out <= 12'h088;
      20'h0a111: out <= 12'h088;
      20'h0a112: out <= 12'h088;
      20'h0a113: out <= 12'h088;
      20'h0a114: out <= 12'h088;
      20'h0a115: out <= 12'h088;
      20'h0a116: out <= 12'h088;
      20'h0a117: out <= 12'h088;
      20'h0a118: out <= 12'h088;
      20'h0a119: out <= 12'h088;
      20'h0a11a: out <= 12'h088;
      20'h0a11b: out <= 12'h088;
      20'h0a11c: out <= 12'h088;
      20'h0a11d: out <= 12'h088;
      20'h0a11e: out <= 12'h088;
      20'h0a11f: out <= 12'h088;
      20'h0a120: out <= 12'h088;
      20'h0a121: out <= 12'h088;
      20'h0a122: out <= 12'h088;
      20'h0a123: out <= 12'h088;
      20'h0a124: out <= 12'h088;
      20'h0a125: out <= 12'h088;
      20'h0a126: out <= 12'h088;
      20'h0a127: out <= 12'h088;
      20'h0a128: out <= 12'h088;
      20'h0a129: out <= 12'h088;
      20'h0a12a: out <= 12'h088;
      20'h0a12b: out <= 12'h088;
      20'h0a12c: out <= 12'h088;
      20'h0a12d: out <= 12'h088;
      20'h0a12e: out <= 12'h088;
      20'h0a12f: out <= 12'h088;
      20'h0a130: out <= 12'h088;
      20'h0a131: out <= 12'h660;
      20'h0a132: out <= 12'h660;
      20'h0a133: out <= 12'h660;
      20'h0a134: out <= 12'h660;
      20'h0a135: out <= 12'h660;
      20'h0a136: out <= 12'h660;
      20'h0a137: out <= 12'h660;
      20'h0a138: out <= 12'h222;
      20'h0a139: out <= 12'h660;
      20'h0a13a: out <= 12'h660;
      20'h0a13b: out <= 12'h660;
      20'h0a13c: out <= 12'hee9;
      20'h0a13d: out <= 12'h660;
      20'h0a13e: out <= 12'h660;
      20'h0a13f: out <= 12'h660;
      20'h0a140: out <= 12'h660;
      20'h0a141: out <= 12'h660;
      20'h0a142: out <= 12'h660;
      20'h0a143: out <= 12'h660;
      20'h0a144: out <= 12'h660;
      20'h0a145: out <= 12'h660;
      20'h0a146: out <= 12'hee9;
      20'h0a147: out <= 12'h660;
      20'h0a148: out <= 12'h603;
      20'h0a149: out <= 12'h603;
      20'h0a14a: out <= 12'h603;
      20'h0a14b: out <= 12'h603;
      20'h0a14c: out <= 12'h4cd;
      20'h0a14d: out <= 12'h4cd;
      20'h0a14e: out <= 12'h000;
      20'h0a14f: out <= 12'h4cd;
      20'h0a150: out <= 12'h000;
      20'h0a151: out <= 12'h4cd;
      20'h0a152: out <= 12'h4cd;
      20'h0a153: out <= 12'h000;
      20'h0a154: out <= 12'h000;
      20'h0a155: out <= 12'h000;
      20'h0a156: out <= 12'h000;
      20'h0a157: out <= 12'h4cd;
      20'h0a158: out <= 12'h4cd;
      20'h0a159: out <= 12'h000;
      20'h0a15a: out <= 12'h000;
      20'h0a15b: out <= 12'h000;
      20'h0a15c: out <= 12'h000;
      20'h0a15d: out <= 12'h000;
      20'h0a15e: out <= 12'h000;
      20'h0a15f: out <= 12'h4cd;
      20'h0a160: out <= 12'h4cd;
      20'h0a161: out <= 12'h4cd;
      20'h0a162: out <= 12'h000;
      20'h0a163: out <= 12'h000;
      20'h0a164: out <= 12'h000;
      20'h0a165: out <= 12'h000;
      20'h0a166: out <= 12'h4cd;
      20'h0a167: out <= 12'h4cd;
      20'h0a168: out <= 12'h4cd;
      20'h0a169: out <= 12'h4cd;
      20'h0a16a: out <= 12'h000;
      20'h0a16b: out <= 12'h000;
      20'h0a16c: out <= 12'h4cd;
      20'h0a16d: out <= 12'h4cd;
      20'h0a16e: out <= 12'h000;
      20'h0a16f: out <= 12'h000;
      20'h0a170: out <= 12'h4cd;
      20'h0a171: out <= 12'h4cd;
      20'h0a172: out <= 12'h000;
      20'h0a173: out <= 12'h000;
      20'h0a174: out <= 12'h000;
      20'h0a175: out <= 12'h000;
      20'h0a176: out <= 12'h000;
      20'h0a177: out <= 12'h000;
      20'h0a178: out <= 12'h000;
      20'h0a179: out <= 12'h4cd;
      20'h0a17a: out <= 12'h4cd;
      20'h0a17b: out <= 12'h000;
      20'h0a17c: out <= 12'h4cd;
      20'h0a17d: out <= 12'h4cd;
      20'h0a17e: out <= 12'h4cd;
      20'h0a17f: out <= 12'h4cd;
      20'h0a180: out <= 12'h4cd;
      20'h0a181: out <= 12'h4cd;
      20'h0a182: out <= 12'h000;
      20'h0a183: out <= 12'h000;
      20'h0a184: out <= 12'h000;
      20'h0a185: out <= 12'h000;
      20'h0a186: out <= 12'h000;
      20'h0a187: out <= 12'h4cd;
      20'h0a188: out <= 12'h4cd;
      20'h0a189: out <= 12'h000;
      20'h0a18a: out <= 12'h000;
      20'h0a18b: out <= 12'h000;
      20'h0a18c: out <= 12'h000;
      20'h0a18d: out <= 12'h4cd;
      20'h0a18e: out <= 12'h4cd;
      20'h0a18f: out <= 12'h4cd;
      20'h0a190: out <= 12'h4cd;
      20'h0a191: out <= 12'h4cd;
      20'h0a192: out <= 12'h000;
      20'h0a193: out <= 12'h000;
      20'h0a194: out <= 12'h000;
      20'h0a195: out <= 12'h4cd;
      20'h0a196: out <= 12'h4cd;
      20'h0a197: out <= 12'h4cd;
      20'h0a198: out <= 12'h4cd;
      20'h0a199: out <= 12'h4cd;
      20'h0a19a: out <= 12'h4cd;
      20'h0a19b: out <= 12'h000;
      20'h0a19c: out <= 12'h603;
      20'h0a19d: out <= 12'h603;
      20'h0a19e: out <= 12'h603;
      20'h0a19f: out <= 12'h603;
      20'h0a1a0: out <= 12'hee9;
      20'h0a1a1: out <= 12'hf87;
      20'h0a1a2: out <= 12'hee9;
      20'h0a1a3: out <= 12'hf87;
      20'h0a1a4: out <= 12'hf87;
      20'h0a1a5: out <= 12'hb27;
      20'h0a1a6: out <= 12'hf87;
      20'h0a1a7: out <= 12'hb27;
      20'h0a1a8: out <= 12'h000;
      20'h0a1a9: out <= 12'h000;
      20'h0a1aa: out <= 12'h000;
      20'h0a1ab: out <= 12'h000;
      20'h0a1ac: out <= 12'h000;
      20'h0a1ad: out <= 12'h000;
      20'h0a1ae: out <= 12'h000;
      20'h0a1af: out <= 12'h000;
      20'h0a1b0: out <= 12'h000;
      20'h0a1b1: out <= 12'hc7f;
      20'h0a1b2: out <= 12'h72f;
      20'h0a1b3: out <= 12'h72f;
      20'h0a1b4: out <= 12'hfff;
      20'h0a1b5: out <= 12'hc7f;
      20'h0a1b6: out <= 12'hc7f;
      20'h0a1b7: out <= 12'h72f;
      20'h0a1b8: out <= 12'h72f;
      20'h0a1b9: out <= 12'h72f;
      20'h0a1ba: out <= 12'hc7f;
      20'h0a1bb: out <= 12'hc7f;
      20'h0a1bc: out <= 12'hfff;
      20'h0a1bd: out <= 12'h72f;
      20'h0a1be: out <= 12'h72f;
      20'h0a1bf: out <= 12'hc7f;
      20'h0a1c0: out <= 12'h000;
      20'h0a1c1: out <= 12'h000;
      20'h0a1c2: out <= 12'h000;
      20'h0a1c3: out <= 12'h000;
      20'h0a1c4: out <= 12'h4cd;
      20'h0a1c5: out <= 12'h000;
      20'h0a1c6: out <= 12'h000;
      20'h0a1c7: out <= 12'h000;
      20'h0a1c8: out <= 12'h4cd;
      20'h0a1c9: out <= 12'h4cd;
      20'h0a1ca: out <= 12'h4cd;
      20'h0a1cb: out <= 12'h4cd;
      20'h0a1cc: out <= 12'h4cd;
      20'h0a1cd: out <= 12'h4cd;
      20'h0a1ce: out <= 12'h4cd;
      20'h0a1cf: out <= 12'h4cd;
      20'h0a1d0: out <= 12'h5ef;
      20'h0a1d1: out <= 12'h5ef;
      20'h0a1d2: out <= 12'h5ef;
      20'h0a1d3: out <= 12'h5ef;
      20'h0a1d4: out <= 12'h5ef;
      20'h0a1d5: out <= 12'h5ef;
      20'h0a1d6: out <= 12'h5ef;
      20'h0a1d7: out <= 12'h5ef;
      20'h0a1d8: out <= 12'h000;
      20'h0a1d9: out <= 12'h000;
      20'h0a1da: out <= 12'h000;
      20'h0a1db: out <= 12'h000;
      20'h0a1dc: out <= 12'h000;
      20'h0a1dd: out <= 12'h000;
      20'h0a1de: out <= 12'h000;
      20'h0a1df: out <= 12'h000;
      20'h0a1e0: out <= 12'h088;
      20'h0a1e1: out <= 12'h088;
      20'h0a1e2: out <= 12'h088;
      20'h0a1e3: out <= 12'h088;
      20'h0a1e4: out <= 12'h088;
      20'h0a1e5: out <= 12'h088;
      20'h0a1e6: out <= 12'h088;
      20'h0a1e7: out <= 12'h088;
      20'h0a1e8: out <= 12'h088;
      20'h0a1e9: out <= 12'h088;
      20'h0a1ea: out <= 12'h088;
      20'h0a1eb: out <= 12'h088;
      20'h0a1ec: out <= 12'h088;
      20'h0a1ed: out <= 12'h088;
      20'h0a1ee: out <= 12'h088;
      20'h0a1ef: out <= 12'h088;
      20'h0a1f0: out <= 12'h088;
      20'h0a1f1: out <= 12'h088;
      20'h0a1f2: out <= 12'h088;
      20'h0a1f3: out <= 12'h088;
      20'h0a1f4: out <= 12'h088;
      20'h0a1f5: out <= 12'h088;
      20'h0a1f6: out <= 12'h088;
      20'h0a1f7: out <= 12'h088;
      20'h0a1f8: out <= 12'h088;
      20'h0a1f9: out <= 12'h088;
      20'h0a1fa: out <= 12'h088;
      20'h0a1fb: out <= 12'h088;
      20'h0a1fc: out <= 12'h088;
      20'h0a1fd: out <= 12'h088;
      20'h0a1fe: out <= 12'h088;
      20'h0a1ff: out <= 12'h088;
      20'h0a200: out <= 12'h088;
      20'h0a201: out <= 12'h088;
      20'h0a202: out <= 12'h088;
      20'h0a203: out <= 12'h088;
      20'h0a204: out <= 12'h088;
      20'h0a205: out <= 12'h088;
      20'h0a206: out <= 12'h088;
      20'h0a207: out <= 12'h088;
      20'h0a208: out <= 12'h088;
      20'h0a209: out <= 12'h088;
      20'h0a20a: out <= 12'h088;
      20'h0a20b: out <= 12'h088;
      20'h0a20c: out <= 12'h088;
      20'h0a20d: out <= 12'h088;
      20'h0a20e: out <= 12'h088;
      20'h0a20f: out <= 12'h088;
      20'h0a210: out <= 12'h088;
      20'h0a211: out <= 12'h088;
      20'h0a212: out <= 12'h088;
      20'h0a213: out <= 12'h088;
      20'h0a214: out <= 12'h088;
      20'h0a215: out <= 12'h088;
      20'h0a216: out <= 12'h088;
      20'h0a217: out <= 12'h088;
      20'h0a218: out <= 12'h088;
      20'h0a219: out <= 12'h088;
      20'h0a21a: out <= 12'h088;
      20'h0a21b: out <= 12'h088;
      20'h0a21c: out <= 12'h088;
      20'h0a21d: out <= 12'h088;
      20'h0a21e: out <= 12'h088;
      20'h0a21f: out <= 12'h088;
      20'h0a220: out <= 12'h088;
      20'h0a221: out <= 12'h088;
      20'h0a222: out <= 12'h088;
      20'h0a223: out <= 12'h088;
      20'h0a224: out <= 12'h088;
      20'h0a225: out <= 12'h088;
      20'h0a226: out <= 12'h088;
      20'h0a227: out <= 12'h088;
      20'h0a228: out <= 12'h088;
      20'h0a229: out <= 12'h088;
      20'h0a22a: out <= 12'h088;
      20'h0a22b: out <= 12'h088;
      20'h0a22c: out <= 12'h088;
      20'h0a22d: out <= 12'h088;
      20'h0a22e: out <= 12'h088;
      20'h0a22f: out <= 12'h088;
      20'h0a230: out <= 12'h088;
      20'h0a231: out <= 12'h088;
      20'h0a232: out <= 12'h088;
      20'h0a233: out <= 12'h088;
      20'h0a234: out <= 12'h088;
      20'h0a235: out <= 12'h088;
      20'h0a236: out <= 12'h088;
      20'h0a237: out <= 12'h088;
      20'h0a238: out <= 12'h088;
      20'h0a239: out <= 12'h088;
      20'h0a23a: out <= 12'h088;
      20'h0a23b: out <= 12'h088;
      20'h0a23c: out <= 12'h088;
      20'h0a23d: out <= 12'h088;
      20'h0a23e: out <= 12'h088;
      20'h0a23f: out <= 12'h088;
      20'h0a240: out <= 12'h088;
      20'h0a241: out <= 12'h088;
      20'h0a242: out <= 12'h088;
      20'h0a243: out <= 12'h088;
      20'h0a244: out <= 12'h088;
      20'h0a245: out <= 12'h088;
      20'h0a246: out <= 12'h088;
      20'h0a247: out <= 12'h088;
      20'h0a248: out <= 12'h088;
      20'h0a249: out <= 12'hbb0;
      20'h0a24a: out <= 12'hbb0;
      20'h0a24b: out <= 12'h660;
      20'h0a24c: out <= 12'h660;
      20'h0a24d: out <= 12'h660;
      20'h0a24e: out <= 12'hee9;
      20'h0a24f: out <= 12'h660;
      20'h0a250: out <= 12'h222;
      20'h0a251: out <= 12'h660;
      20'h0a252: out <= 12'hee9;
      20'h0a253: out <= 12'h660;
      20'h0a254: out <= 12'hee9;
      20'h0a255: out <= 12'h660;
      20'h0a256: out <= 12'hbb0;
      20'h0a257: out <= 12'hbb0;
      20'h0a258: out <= 12'hbb0;
      20'h0a259: out <= 12'hbb0;
      20'h0a25a: out <= 12'hbb0;
      20'h0a25b: out <= 12'h660;
      20'h0a25c: out <= 12'h660;
      20'h0a25d: out <= 12'h660;
      20'h0a25e: out <= 12'h660;
      20'h0a25f: out <= 12'h660;
      20'h0a260: out <= 12'h603;
      20'h0a261: out <= 12'h603;
      20'h0a262: out <= 12'h603;
      20'h0a263: out <= 12'h603;
      20'h0a264: out <= 12'h4cd;
      20'h0a265: out <= 12'h4cd;
      20'h0a266: out <= 12'h4cd;
      20'h0a267: out <= 12'h000;
      20'h0a268: out <= 12'h000;
      20'h0a269: out <= 12'h4cd;
      20'h0a26a: out <= 12'h4cd;
      20'h0a26b: out <= 12'h000;
      20'h0a26c: out <= 12'h000;
      20'h0a26d: out <= 12'h000;
      20'h0a26e: out <= 12'h000;
      20'h0a26f: out <= 12'h4cd;
      20'h0a270: out <= 12'h4cd;
      20'h0a271: out <= 12'h000;
      20'h0a272: out <= 12'h000;
      20'h0a273: out <= 12'h000;
      20'h0a274: out <= 12'h000;
      20'h0a275: out <= 12'h4cd;
      20'h0a276: out <= 12'h4cd;
      20'h0a277: out <= 12'h4cd;
      20'h0a278: out <= 12'h000;
      20'h0a279: out <= 12'h000;
      20'h0a27a: out <= 12'h000;
      20'h0a27b: out <= 12'h000;
      20'h0a27c: out <= 12'h000;
      20'h0a27d: out <= 12'h000;
      20'h0a27e: out <= 12'h000;
      20'h0a27f: out <= 12'h000;
      20'h0a280: out <= 12'h000;
      20'h0a281: out <= 12'h4cd;
      20'h0a282: out <= 12'h4cd;
      20'h0a283: out <= 12'h000;
      20'h0a284: out <= 12'h4cd;
      20'h0a285: out <= 12'h4cd;
      20'h0a286: out <= 12'h4cd;
      20'h0a287: out <= 12'h4cd;
      20'h0a288: out <= 12'h4cd;
      20'h0a289: out <= 12'h4cd;
      20'h0a28a: out <= 12'h4cd;
      20'h0a28b: out <= 12'h000;
      20'h0a28c: out <= 12'h000;
      20'h0a28d: out <= 12'h000;
      20'h0a28e: out <= 12'h000;
      20'h0a28f: out <= 12'h000;
      20'h0a290: out <= 12'h000;
      20'h0a291: out <= 12'h4cd;
      20'h0a292: out <= 12'h4cd;
      20'h0a293: out <= 12'h000;
      20'h0a294: out <= 12'h4cd;
      20'h0a295: out <= 12'h4cd;
      20'h0a296: out <= 12'h000;
      20'h0a297: out <= 12'h000;
      20'h0a298: out <= 12'h000;
      20'h0a299: out <= 12'h4cd;
      20'h0a29a: out <= 12'h4cd;
      20'h0a29b: out <= 12'h000;
      20'h0a29c: out <= 12'h000;
      20'h0a29d: out <= 12'h000;
      20'h0a29e: out <= 12'h4cd;
      20'h0a29f: out <= 12'h4cd;
      20'h0a2a0: out <= 12'h000;
      20'h0a2a1: out <= 12'h000;
      20'h0a2a2: out <= 12'h000;
      20'h0a2a3: out <= 12'h000;
      20'h0a2a4: out <= 12'h4cd;
      20'h0a2a5: out <= 12'h4cd;
      20'h0a2a6: out <= 12'h000;
      20'h0a2a7: out <= 12'h000;
      20'h0a2a8: out <= 12'h000;
      20'h0a2a9: out <= 12'h4cd;
      20'h0a2aa: out <= 12'h4cd;
      20'h0a2ab: out <= 12'h000;
      20'h0a2ac: out <= 12'h000;
      20'h0a2ad: out <= 12'h000;
      20'h0a2ae: out <= 12'h000;
      20'h0a2af: out <= 12'h000;
      20'h0a2b0: out <= 12'h000;
      20'h0a2b1: out <= 12'h4cd;
      20'h0a2b2: out <= 12'h4cd;
      20'h0a2b3: out <= 12'h000;
      20'h0a2b4: out <= 12'h603;
      20'h0a2b5: out <= 12'h603;
      20'h0a2b6: out <= 12'h603;
      20'h0a2b7: out <= 12'h603;
      20'h0a2b8: out <= 12'hee9;
      20'h0a2b9: out <= 12'hf87;
      20'h0a2ba: out <= 12'hee9;
      20'h0a2bb: out <= 12'hf87;
      20'h0a2bc: out <= 12'hf87;
      20'h0a2bd: out <= 12'hb27;
      20'h0a2be: out <= 12'hf87;
      20'h0a2bf: out <= 12'hb27;
      20'h0a2c0: out <= 12'h000;
      20'h0a2c1: out <= 12'h000;
      20'h0a2c2: out <= 12'h000;
      20'h0a2c3: out <= 12'h000;
      20'h0a2c4: out <= 12'h000;
      20'h0a2c5: out <= 12'h000;
      20'h0a2c6: out <= 12'h000;
      20'h0a2c7: out <= 12'h000;
      20'h0a2c8: out <= 12'h000;
      20'h0a2c9: out <= 12'hc7f;
      20'h0a2ca: out <= 12'hfff;
      20'h0a2cb: out <= 12'hc7f;
      20'h0a2cc: out <= 12'h72f;
      20'h0a2cd: out <= 12'hfff;
      20'h0a2ce: out <= 12'hc7f;
      20'h0a2cf: out <= 12'hc7f;
      20'h0a2d0: out <= 12'hc7f;
      20'h0a2d1: out <= 12'hc7f;
      20'h0a2d2: out <= 12'hc7f;
      20'h0a2d3: out <= 12'hfff;
      20'h0a2d4: out <= 12'h72f;
      20'h0a2d5: out <= 12'hc7f;
      20'h0a2d6: out <= 12'hfff;
      20'h0a2d7: out <= 12'hc7f;
      20'h0a2d8: out <= 12'h000;
      20'h0a2d9: out <= 12'h000;
      20'h0a2da: out <= 12'h000;
      20'h0a2db: out <= 12'h4cd;
      20'h0a2dc: out <= 12'h000;
      20'h0a2dd: out <= 12'h4cd;
      20'h0a2de: out <= 12'h000;
      20'h0a2df: out <= 12'h000;
      20'h0a2e0: out <= 12'h4cd;
      20'h0a2e1: out <= 12'h4cd;
      20'h0a2e2: out <= 12'h4cd;
      20'h0a2e3: out <= 12'h4cd;
      20'h0a2e4: out <= 12'h4cd;
      20'h0a2e5: out <= 12'h4cd;
      20'h0a2e6: out <= 12'h4cd;
      20'h0a2e7: out <= 12'h4cd;
      20'h0a2e8: out <= 12'h5ef;
      20'h0a2e9: out <= 12'h5ef;
      20'h0a2ea: out <= 12'h5ef;
      20'h0a2eb: out <= 12'h5ef;
      20'h0a2ec: out <= 12'h5ef;
      20'h0a2ed: out <= 12'h5ef;
      20'h0a2ee: out <= 12'h5ef;
      20'h0a2ef: out <= 12'h5ef;
      20'h0a2f0: out <= 12'h000;
      20'h0a2f1: out <= 12'h000;
      20'h0a2f2: out <= 12'h000;
      20'h0a2f3: out <= 12'h000;
      20'h0a2f4: out <= 12'h000;
      20'h0a2f5: out <= 12'h000;
      20'h0a2f6: out <= 12'h000;
      20'h0a2f7: out <= 12'h000;
      20'h0a2f8: out <= 12'h088;
      20'h0a2f9: out <= 12'h088;
      20'h0a2fa: out <= 12'h088;
      20'h0a2fb: out <= 12'h088;
      20'h0a2fc: out <= 12'h088;
      20'h0a2fd: out <= 12'h088;
      20'h0a2fe: out <= 12'h088;
      20'h0a2ff: out <= 12'h088;
      20'h0a300: out <= 12'h088;
      20'h0a301: out <= 12'h088;
      20'h0a302: out <= 12'h088;
      20'h0a303: out <= 12'h088;
      20'h0a304: out <= 12'h088;
      20'h0a305: out <= 12'h088;
      20'h0a306: out <= 12'h088;
      20'h0a307: out <= 12'h088;
      20'h0a308: out <= 12'h088;
      20'h0a309: out <= 12'h088;
      20'h0a30a: out <= 12'h088;
      20'h0a30b: out <= 12'h088;
      20'h0a30c: out <= 12'h088;
      20'h0a30d: out <= 12'h088;
      20'h0a30e: out <= 12'h088;
      20'h0a30f: out <= 12'h088;
      20'h0a310: out <= 12'h088;
      20'h0a311: out <= 12'h088;
      20'h0a312: out <= 12'h088;
      20'h0a313: out <= 12'h088;
      20'h0a314: out <= 12'h088;
      20'h0a315: out <= 12'h088;
      20'h0a316: out <= 12'h088;
      20'h0a317: out <= 12'h088;
      20'h0a318: out <= 12'h088;
      20'h0a319: out <= 12'h088;
      20'h0a31a: out <= 12'h088;
      20'h0a31b: out <= 12'h088;
      20'h0a31c: out <= 12'h088;
      20'h0a31d: out <= 12'h088;
      20'h0a31e: out <= 12'h088;
      20'h0a31f: out <= 12'h088;
      20'h0a320: out <= 12'h088;
      20'h0a321: out <= 12'h088;
      20'h0a322: out <= 12'h088;
      20'h0a323: out <= 12'h088;
      20'h0a324: out <= 12'h088;
      20'h0a325: out <= 12'h088;
      20'h0a326: out <= 12'h088;
      20'h0a327: out <= 12'h088;
      20'h0a328: out <= 12'h088;
      20'h0a329: out <= 12'h088;
      20'h0a32a: out <= 12'h088;
      20'h0a32b: out <= 12'h088;
      20'h0a32c: out <= 12'h088;
      20'h0a32d: out <= 12'h088;
      20'h0a32e: out <= 12'h088;
      20'h0a32f: out <= 12'h088;
      20'h0a330: out <= 12'h088;
      20'h0a331: out <= 12'h088;
      20'h0a332: out <= 12'h088;
      20'h0a333: out <= 12'h088;
      20'h0a334: out <= 12'h088;
      20'h0a335: out <= 12'h088;
      20'h0a336: out <= 12'h088;
      20'h0a337: out <= 12'h088;
      20'h0a338: out <= 12'h088;
      20'h0a339: out <= 12'h088;
      20'h0a33a: out <= 12'h088;
      20'h0a33b: out <= 12'h088;
      20'h0a33c: out <= 12'h088;
      20'h0a33d: out <= 12'h088;
      20'h0a33e: out <= 12'h088;
      20'h0a33f: out <= 12'h088;
      20'h0a340: out <= 12'h088;
      20'h0a341: out <= 12'h088;
      20'h0a342: out <= 12'h088;
      20'h0a343: out <= 12'h088;
      20'h0a344: out <= 12'h088;
      20'h0a345: out <= 12'h088;
      20'h0a346: out <= 12'h088;
      20'h0a347: out <= 12'h088;
      20'h0a348: out <= 12'h088;
      20'h0a349: out <= 12'h088;
      20'h0a34a: out <= 12'h088;
      20'h0a34b: out <= 12'h088;
      20'h0a34c: out <= 12'h088;
      20'h0a34d: out <= 12'h088;
      20'h0a34e: out <= 12'h088;
      20'h0a34f: out <= 12'h088;
      20'h0a350: out <= 12'h088;
      20'h0a351: out <= 12'h088;
      20'h0a352: out <= 12'h088;
      20'h0a353: out <= 12'h088;
      20'h0a354: out <= 12'h088;
      20'h0a355: out <= 12'h088;
      20'h0a356: out <= 12'h088;
      20'h0a357: out <= 12'h088;
      20'h0a358: out <= 12'h088;
      20'h0a359: out <= 12'h088;
      20'h0a35a: out <= 12'h088;
      20'h0a35b: out <= 12'h088;
      20'h0a35c: out <= 12'h088;
      20'h0a35d: out <= 12'h088;
      20'h0a35e: out <= 12'h088;
      20'h0a35f: out <= 12'h088;
      20'h0a360: out <= 12'h088;
      20'h0a361: out <= 12'hee9;
      20'h0a362: out <= 12'hbb0;
      20'h0a363: out <= 12'h660;
      20'h0a364: out <= 12'h660;
      20'h0a365: out <= 12'h660;
      20'h0a366: out <= 12'h660;
      20'h0a367: out <= 12'h660;
      20'h0a368: out <= 12'h222;
      20'h0a369: out <= 12'h660;
      20'h0a36a: out <= 12'h660;
      20'h0a36b: out <= 12'h660;
      20'h0a36c: out <= 12'hee9;
      20'h0a36d: out <= 12'h660;
      20'h0a36e: out <= 12'hbb0;
      20'h0a36f: out <= 12'h660;
      20'h0a370: out <= 12'hee9;
      20'h0a371: out <= 12'hee9;
      20'h0a372: out <= 12'hbb0;
      20'h0a373: out <= 12'h660;
      20'h0a374: out <= 12'h660;
      20'h0a375: out <= 12'h660;
      20'h0a376: out <= 12'hee9;
      20'h0a377: out <= 12'h660;
      20'h0a378: out <= 12'h603;
      20'h0a379: out <= 12'h603;
      20'h0a37a: out <= 12'h603;
      20'h0a37b: out <= 12'h603;
      20'h0a37c: out <= 12'h4cd;
      20'h0a37d: out <= 12'h4cd;
      20'h0a37e: out <= 12'h000;
      20'h0a37f: out <= 12'h000;
      20'h0a380: out <= 12'h000;
      20'h0a381: out <= 12'h4cd;
      20'h0a382: out <= 12'h4cd;
      20'h0a383: out <= 12'h000;
      20'h0a384: out <= 12'h000;
      20'h0a385: out <= 12'h000;
      20'h0a386: out <= 12'h000;
      20'h0a387: out <= 12'h4cd;
      20'h0a388: out <= 12'h4cd;
      20'h0a389: out <= 12'h000;
      20'h0a38a: out <= 12'h000;
      20'h0a38b: out <= 12'h000;
      20'h0a38c: out <= 12'h4cd;
      20'h0a38d: out <= 12'h4cd;
      20'h0a38e: out <= 12'h000;
      20'h0a38f: out <= 12'h000;
      20'h0a390: out <= 12'h000;
      20'h0a391: out <= 12'h000;
      20'h0a392: out <= 12'h000;
      20'h0a393: out <= 12'h000;
      20'h0a394: out <= 12'h4cd;
      20'h0a395: out <= 12'h4cd;
      20'h0a396: out <= 12'h000;
      20'h0a397: out <= 12'h000;
      20'h0a398: out <= 12'h000;
      20'h0a399: out <= 12'h4cd;
      20'h0a39a: out <= 12'h4cd;
      20'h0a39b: out <= 12'h000;
      20'h0a39c: out <= 12'h000;
      20'h0a39d: out <= 12'h000;
      20'h0a39e: out <= 12'h000;
      20'h0a39f: out <= 12'h000;
      20'h0a3a0: out <= 12'h4cd;
      20'h0a3a1: out <= 12'h4cd;
      20'h0a3a2: out <= 12'h000;
      20'h0a3a3: out <= 12'h000;
      20'h0a3a4: out <= 12'h4cd;
      20'h0a3a5: out <= 12'h4cd;
      20'h0a3a6: out <= 12'h000;
      20'h0a3a7: out <= 12'h000;
      20'h0a3a8: out <= 12'h000;
      20'h0a3a9: out <= 12'h4cd;
      20'h0a3aa: out <= 12'h4cd;
      20'h0a3ab: out <= 12'h000;
      20'h0a3ac: out <= 12'h4cd;
      20'h0a3ad: out <= 12'h4cd;
      20'h0a3ae: out <= 12'h000;
      20'h0a3af: out <= 12'h000;
      20'h0a3b0: out <= 12'h000;
      20'h0a3b1: out <= 12'h4cd;
      20'h0a3b2: out <= 12'h4cd;
      20'h0a3b3: out <= 12'h000;
      20'h0a3b4: out <= 12'h000;
      20'h0a3b5: out <= 12'h000;
      20'h0a3b6: out <= 12'h4cd;
      20'h0a3b7: out <= 12'h4cd;
      20'h0a3b8: out <= 12'h000;
      20'h0a3b9: out <= 12'h000;
      20'h0a3ba: out <= 12'h000;
      20'h0a3bb: out <= 12'h000;
      20'h0a3bc: out <= 12'h4cd;
      20'h0a3bd: out <= 12'h4cd;
      20'h0a3be: out <= 12'h000;
      20'h0a3bf: out <= 12'h000;
      20'h0a3c0: out <= 12'h000;
      20'h0a3c1: out <= 12'h4cd;
      20'h0a3c2: out <= 12'h4cd;
      20'h0a3c3: out <= 12'h000;
      20'h0a3c4: out <= 12'h000;
      20'h0a3c5: out <= 12'h000;
      20'h0a3c6: out <= 12'h000;
      20'h0a3c7: out <= 12'h000;
      20'h0a3c8: out <= 12'h4cd;
      20'h0a3c9: out <= 12'h4cd;
      20'h0a3ca: out <= 12'h000;
      20'h0a3cb: out <= 12'h000;
      20'h0a3cc: out <= 12'h603;
      20'h0a3cd: out <= 12'h603;
      20'h0a3ce: out <= 12'h603;
      20'h0a3cf: out <= 12'h603;
      20'h0a3d0: out <= 12'hee9;
      20'h0a3d1: out <= 12'hf87;
      20'h0a3d2: out <= 12'hee9;
      20'h0a3d3: out <= 12'hb27;
      20'h0a3d4: out <= 12'hb27;
      20'h0a3d5: out <= 12'hb27;
      20'h0a3d6: out <= 12'hf87;
      20'h0a3d7: out <= 12'hb27;
      20'h0a3d8: out <= 12'h000;
      20'h0a3d9: out <= 12'h000;
      20'h0a3da: out <= 12'h000;
      20'h0a3db: out <= 12'h000;
      20'h0a3dc: out <= 12'h000;
      20'h0a3dd: out <= 12'h000;
      20'h0a3de: out <= 12'h000;
      20'h0a3df: out <= 12'h000;
      20'h0a3e0: out <= 12'h000;
      20'h0a3e1: out <= 12'hc7f;
      20'h0a3e2: out <= 12'h72f;
      20'h0a3e3: out <= 12'hc7f;
      20'h0a3e4: out <= 12'h000;
      20'h0a3e5: out <= 12'h72f;
      20'h0a3e6: out <= 12'h72f;
      20'h0a3e7: out <= 12'h72f;
      20'h0a3e8: out <= 12'h72f;
      20'h0a3e9: out <= 12'h72f;
      20'h0a3ea: out <= 12'h72f;
      20'h0a3eb: out <= 12'h72f;
      20'h0a3ec: out <= 12'h000;
      20'h0a3ed: out <= 12'hc7f;
      20'h0a3ee: out <= 12'h72f;
      20'h0a3ef: out <= 12'hc7f;
      20'h0a3f0: out <= 12'h000;
      20'h0a3f1: out <= 12'h000;
      20'h0a3f2: out <= 12'h4cd;
      20'h0a3f3: out <= 12'h000;
      20'h0a3f4: out <= 12'h000;
      20'h0a3f5: out <= 12'h000;
      20'h0a3f6: out <= 12'h4cd;
      20'h0a3f7: out <= 12'h000;
      20'h0a3f8: out <= 12'h4cd;
      20'h0a3f9: out <= 12'h4cd;
      20'h0a3fa: out <= 12'h4cd;
      20'h0a3fb: out <= 12'h4cd;
      20'h0a3fc: out <= 12'h4cd;
      20'h0a3fd: out <= 12'h4cd;
      20'h0a3fe: out <= 12'h4cd;
      20'h0a3ff: out <= 12'h4cd;
      20'h0a400: out <= 12'h5ef;
      20'h0a401: out <= 12'h5ef;
      20'h0a402: out <= 12'h5ef;
      20'h0a403: out <= 12'h5ef;
      20'h0a404: out <= 12'h5ef;
      20'h0a405: out <= 12'h5ef;
      20'h0a406: out <= 12'h5ef;
      20'h0a407: out <= 12'h5ef;
      20'h0a408: out <= 12'h000;
      20'h0a409: out <= 12'h000;
      20'h0a40a: out <= 12'h000;
      20'h0a40b: out <= 12'h000;
      20'h0a40c: out <= 12'h000;
      20'h0a40d: out <= 12'h000;
      20'h0a40e: out <= 12'h000;
      20'h0a40f: out <= 12'h000;
      20'h0a410: out <= 12'h088;
      20'h0a411: out <= 12'h088;
      20'h0a412: out <= 12'h088;
      20'h0a413: out <= 12'h088;
      20'h0a414: out <= 12'h088;
      20'h0a415: out <= 12'h088;
      20'h0a416: out <= 12'h088;
      20'h0a417: out <= 12'h088;
      20'h0a418: out <= 12'h088;
      20'h0a419: out <= 12'h088;
      20'h0a41a: out <= 12'h088;
      20'h0a41b: out <= 12'h088;
      20'h0a41c: out <= 12'h088;
      20'h0a41d: out <= 12'h088;
      20'h0a41e: out <= 12'h088;
      20'h0a41f: out <= 12'h088;
      20'h0a420: out <= 12'h088;
      20'h0a421: out <= 12'h088;
      20'h0a422: out <= 12'h088;
      20'h0a423: out <= 12'h088;
      20'h0a424: out <= 12'h088;
      20'h0a425: out <= 12'h088;
      20'h0a426: out <= 12'h088;
      20'h0a427: out <= 12'h088;
      20'h0a428: out <= 12'h088;
      20'h0a429: out <= 12'h088;
      20'h0a42a: out <= 12'h088;
      20'h0a42b: out <= 12'h088;
      20'h0a42c: out <= 12'h088;
      20'h0a42d: out <= 12'h088;
      20'h0a42e: out <= 12'h088;
      20'h0a42f: out <= 12'h088;
      20'h0a430: out <= 12'h088;
      20'h0a431: out <= 12'h088;
      20'h0a432: out <= 12'h088;
      20'h0a433: out <= 12'h088;
      20'h0a434: out <= 12'h088;
      20'h0a435: out <= 12'h088;
      20'h0a436: out <= 12'h088;
      20'h0a437: out <= 12'h088;
      20'h0a438: out <= 12'h088;
      20'h0a439: out <= 12'h088;
      20'h0a43a: out <= 12'h088;
      20'h0a43b: out <= 12'h088;
      20'h0a43c: out <= 12'h088;
      20'h0a43d: out <= 12'h088;
      20'h0a43e: out <= 12'h088;
      20'h0a43f: out <= 12'h088;
      20'h0a440: out <= 12'h088;
      20'h0a441: out <= 12'h088;
      20'h0a442: out <= 12'h088;
      20'h0a443: out <= 12'h088;
      20'h0a444: out <= 12'h088;
      20'h0a445: out <= 12'h088;
      20'h0a446: out <= 12'h088;
      20'h0a447: out <= 12'h088;
      20'h0a448: out <= 12'h088;
      20'h0a449: out <= 12'h088;
      20'h0a44a: out <= 12'h088;
      20'h0a44b: out <= 12'h088;
      20'h0a44c: out <= 12'h088;
      20'h0a44d: out <= 12'h088;
      20'h0a44e: out <= 12'h088;
      20'h0a44f: out <= 12'h088;
      20'h0a450: out <= 12'h088;
      20'h0a451: out <= 12'h088;
      20'h0a452: out <= 12'h088;
      20'h0a453: out <= 12'h088;
      20'h0a454: out <= 12'h088;
      20'h0a455: out <= 12'h088;
      20'h0a456: out <= 12'h088;
      20'h0a457: out <= 12'h088;
      20'h0a458: out <= 12'h088;
      20'h0a459: out <= 12'h088;
      20'h0a45a: out <= 12'h088;
      20'h0a45b: out <= 12'h088;
      20'h0a45c: out <= 12'h088;
      20'h0a45d: out <= 12'h088;
      20'h0a45e: out <= 12'h088;
      20'h0a45f: out <= 12'h088;
      20'h0a460: out <= 12'h088;
      20'h0a461: out <= 12'h088;
      20'h0a462: out <= 12'h088;
      20'h0a463: out <= 12'h088;
      20'h0a464: out <= 12'h088;
      20'h0a465: out <= 12'h088;
      20'h0a466: out <= 12'h088;
      20'h0a467: out <= 12'h088;
      20'h0a468: out <= 12'h088;
      20'h0a469: out <= 12'h088;
      20'h0a46a: out <= 12'h088;
      20'h0a46b: out <= 12'h088;
      20'h0a46c: out <= 12'h088;
      20'h0a46d: out <= 12'h088;
      20'h0a46e: out <= 12'h088;
      20'h0a46f: out <= 12'h088;
      20'h0a470: out <= 12'h088;
      20'h0a471: out <= 12'h088;
      20'h0a472: out <= 12'h088;
      20'h0a473: out <= 12'h088;
      20'h0a474: out <= 12'h088;
      20'h0a475: out <= 12'h088;
      20'h0a476: out <= 12'h088;
      20'h0a477: out <= 12'h088;
      20'h0a478: out <= 12'h088;
      20'h0a479: out <= 12'hee9;
      20'h0a47a: out <= 12'hbb0;
      20'h0a47b: out <= 12'h660;
      20'h0a47c: out <= 12'h660;
      20'h0a47d: out <= 12'h660;
      20'h0a47e: out <= 12'hee9;
      20'h0a47f: out <= 12'h660;
      20'h0a480: out <= 12'h222;
      20'h0a481: out <= 12'h660;
      20'h0a482: out <= 12'hee9;
      20'h0a483: out <= 12'h660;
      20'h0a484: out <= 12'hee9;
      20'h0a485: out <= 12'h660;
      20'h0a486: out <= 12'hbb0;
      20'h0a487: out <= 12'h660;
      20'h0a488: out <= 12'hbb0;
      20'h0a489: out <= 12'hee9;
      20'h0a48a: out <= 12'hbb0;
      20'h0a48b: out <= 12'h660;
      20'h0a48c: out <= 12'h660;
      20'h0a48d: out <= 12'h660;
      20'h0a48e: out <= 12'h660;
      20'h0a48f: out <= 12'h660;
      20'h0a490: out <= 12'h603;
      20'h0a491: out <= 12'h603;
      20'h0a492: out <= 12'h603;
      20'h0a493: out <= 12'h603;
      20'h0a494: out <= 12'h000;
      20'h0a495: out <= 12'h4cd;
      20'h0a496: out <= 12'h4cd;
      20'h0a497: out <= 12'h4cd;
      20'h0a498: out <= 12'h4cd;
      20'h0a499: out <= 12'h4cd;
      20'h0a49a: out <= 12'h000;
      20'h0a49b: out <= 12'h000;
      20'h0a49c: out <= 12'h000;
      20'h0a49d: out <= 12'h000;
      20'h0a49e: out <= 12'h000;
      20'h0a49f: out <= 12'h4cd;
      20'h0a4a0: out <= 12'h4cd;
      20'h0a4a1: out <= 12'h000;
      20'h0a4a2: out <= 12'h000;
      20'h0a4a3: out <= 12'h000;
      20'h0a4a4: out <= 12'h4cd;
      20'h0a4a5: out <= 12'h4cd;
      20'h0a4a6: out <= 12'h4cd;
      20'h0a4a7: out <= 12'h4cd;
      20'h0a4a8: out <= 12'h4cd;
      20'h0a4a9: out <= 12'h4cd;
      20'h0a4aa: out <= 12'h4cd;
      20'h0a4ab: out <= 12'h000;
      20'h0a4ac: out <= 12'h000;
      20'h0a4ad: out <= 12'h4cd;
      20'h0a4ae: out <= 12'h4cd;
      20'h0a4af: out <= 12'h4cd;
      20'h0a4b0: out <= 12'h4cd;
      20'h0a4b1: out <= 12'h4cd;
      20'h0a4b2: out <= 12'h000;
      20'h0a4b3: out <= 12'h000;
      20'h0a4b4: out <= 12'h000;
      20'h0a4b5: out <= 12'h000;
      20'h0a4b6: out <= 12'h000;
      20'h0a4b7: out <= 12'h000;
      20'h0a4b8: out <= 12'h4cd;
      20'h0a4b9: out <= 12'h4cd;
      20'h0a4ba: out <= 12'h000;
      20'h0a4bb: out <= 12'h000;
      20'h0a4bc: out <= 12'h000;
      20'h0a4bd: out <= 12'h4cd;
      20'h0a4be: out <= 12'h4cd;
      20'h0a4bf: out <= 12'h4cd;
      20'h0a4c0: out <= 12'h4cd;
      20'h0a4c1: out <= 12'h4cd;
      20'h0a4c2: out <= 12'h000;
      20'h0a4c3: out <= 12'h000;
      20'h0a4c4: out <= 12'h000;
      20'h0a4c5: out <= 12'h4cd;
      20'h0a4c6: out <= 12'h4cd;
      20'h0a4c7: out <= 12'h4cd;
      20'h0a4c8: out <= 12'h4cd;
      20'h0a4c9: out <= 12'h4cd;
      20'h0a4ca: out <= 12'h000;
      20'h0a4cb: out <= 12'h000;
      20'h0a4cc: out <= 12'h000;
      20'h0a4cd: out <= 12'h000;
      20'h0a4ce: out <= 12'h4cd;
      20'h0a4cf: out <= 12'h4cd;
      20'h0a4d0: out <= 12'h000;
      20'h0a4d1: out <= 12'h000;
      20'h0a4d2: out <= 12'h000;
      20'h0a4d3: out <= 12'h000;
      20'h0a4d4: out <= 12'h000;
      20'h0a4d5: out <= 12'h4cd;
      20'h0a4d6: out <= 12'h4cd;
      20'h0a4d7: out <= 12'h4cd;
      20'h0a4d8: out <= 12'h4cd;
      20'h0a4d9: out <= 12'h4cd;
      20'h0a4da: out <= 12'h000;
      20'h0a4db: out <= 12'h000;
      20'h0a4dc: out <= 12'h000;
      20'h0a4dd: out <= 12'h4cd;
      20'h0a4de: out <= 12'h4cd;
      20'h0a4df: out <= 12'h4cd;
      20'h0a4e0: out <= 12'h4cd;
      20'h0a4e1: out <= 12'h000;
      20'h0a4e2: out <= 12'h000;
      20'h0a4e3: out <= 12'h000;
      20'h0a4e4: out <= 12'h603;
      20'h0a4e5: out <= 12'h603;
      20'h0a4e6: out <= 12'h603;
      20'h0a4e7: out <= 12'h603;
      20'h0a4e8: out <= 12'hee9;
      20'h0a4e9: out <= 12'hf87;
      20'h0a4ea: out <= 12'hf87;
      20'h0a4eb: out <= 12'hf87;
      20'h0a4ec: out <= 12'hf87;
      20'h0a4ed: out <= 12'hf87;
      20'h0a4ee: out <= 12'hf87;
      20'h0a4ef: out <= 12'hb27;
      20'h0a4f0: out <= 12'h000;
      20'h0a4f1: out <= 12'h000;
      20'h0a4f2: out <= 12'h000;
      20'h0a4f3: out <= 12'h000;
      20'h0a4f4: out <= 12'h000;
      20'h0a4f5: out <= 12'h000;
      20'h0a4f6: out <= 12'h000;
      20'h0a4f7: out <= 12'h000;
      20'h0a4f8: out <= 12'h000;
      20'h0a4f9: out <= 12'hc7f;
      20'h0a4fa: out <= 12'hfff;
      20'h0a4fb: out <= 12'hc7f;
      20'h0a4fc: out <= 12'h000;
      20'h0a4fd: out <= 12'h000;
      20'h0a4fe: out <= 12'h000;
      20'h0a4ff: out <= 12'h000;
      20'h0a500: out <= 12'h000;
      20'h0a501: out <= 12'h000;
      20'h0a502: out <= 12'h000;
      20'h0a503: out <= 12'h000;
      20'h0a504: out <= 12'h000;
      20'h0a505: out <= 12'hc7f;
      20'h0a506: out <= 12'hfff;
      20'h0a507: out <= 12'hc7f;
      20'h0a508: out <= 12'h000;
      20'h0a509: out <= 12'h000;
      20'h0a50a: out <= 12'h000;
      20'h0a50b: out <= 12'h000;
      20'h0a50c: out <= 12'h000;
      20'h0a50d: out <= 12'h000;
      20'h0a50e: out <= 12'h000;
      20'h0a50f: out <= 12'h000;
      20'h0a510: out <= 12'h4cd;
      20'h0a511: out <= 12'h4cd;
      20'h0a512: out <= 12'h4cd;
      20'h0a513: out <= 12'h4cd;
      20'h0a514: out <= 12'h4cd;
      20'h0a515: out <= 12'h4cd;
      20'h0a516: out <= 12'h4cd;
      20'h0a517: out <= 12'h4cd;
      20'h0a518: out <= 12'h5ef;
      20'h0a519: out <= 12'h5ef;
      20'h0a51a: out <= 12'h5ef;
      20'h0a51b: out <= 12'h5ef;
      20'h0a51c: out <= 12'h5ef;
      20'h0a51d: out <= 12'h5ef;
      20'h0a51e: out <= 12'h5ef;
      20'h0a51f: out <= 12'h5ef;
      20'h0a520: out <= 12'h000;
      20'h0a521: out <= 12'h000;
      20'h0a522: out <= 12'h000;
      20'h0a523: out <= 12'h000;
      20'h0a524: out <= 12'h000;
      20'h0a525: out <= 12'h000;
      20'h0a526: out <= 12'h000;
      20'h0a527: out <= 12'h000;
      20'h0a528: out <= 12'h088;
      20'h0a529: out <= 12'h088;
      20'h0a52a: out <= 12'h088;
      20'h0a52b: out <= 12'h088;
      20'h0a52c: out <= 12'h088;
      20'h0a52d: out <= 12'h088;
      20'h0a52e: out <= 12'h088;
      20'h0a52f: out <= 12'h088;
      20'h0a530: out <= 12'h088;
      20'h0a531: out <= 12'h088;
      20'h0a532: out <= 12'h088;
      20'h0a533: out <= 12'h088;
      20'h0a534: out <= 12'h088;
      20'h0a535: out <= 12'h088;
      20'h0a536: out <= 12'h088;
      20'h0a537: out <= 12'h088;
      20'h0a538: out <= 12'h088;
      20'h0a539: out <= 12'h088;
      20'h0a53a: out <= 12'h088;
      20'h0a53b: out <= 12'h088;
      20'h0a53c: out <= 12'h088;
      20'h0a53d: out <= 12'h088;
      20'h0a53e: out <= 12'h088;
      20'h0a53f: out <= 12'h088;
      20'h0a540: out <= 12'h088;
      20'h0a541: out <= 12'h088;
      20'h0a542: out <= 12'h088;
      20'h0a543: out <= 12'h088;
      20'h0a544: out <= 12'h088;
      20'h0a545: out <= 12'h088;
      20'h0a546: out <= 12'h088;
      20'h0a547: out <= 12'h088;
      20'h0a548: out <= 12'h088;
      20'h0a549: out <= 12'h088;
      20'h0a54a: out <= 12'h088;
      20'h0a54b: out <= 12'h088;
      20'h0a54c: out <= 12'h088;
      20'h0a54d: out <= 12'h088;
      20'h0a54e: out <= 12'h088;
      20'h0a54f: out <= 12'h088;
      20'h0a550: out <= 12'h088;
      20'h0a551: out <= 12'h088;
      20'h0a552: out <= 12'h088;
      20'h0a553: out <= 12'h088;
      20'h0a554: out <= 12'h088;
      20'h0a555: out <= 12'h088;
      20'h0a556: out <= 12'h088;
      20'h0a557: out <= 12'h088;
      20'h0a558: out <= 12'h088;
      20'h0a559: out <= 12'h088;
      20'h0a55a: out <= 12'h088;
      20'h0a55b: out <= 12'h088;
      20'h0a55c: out <= 12'h088;
      20'h0a55d: out <= 12'h088;
      20'h0a55e: out <= 12'h088;
      20'h0a55f: out <= 12'h088;
      20'h0a560: out <= 12'h088;
      20'h0a561: out <= 12'h088;
      20'h0a562: out <= 12'h088;
      20'h0a563: out <= 12'h088;
      20'h0a564: out <= 12'h088;
      20'h0a565: out <= 12'h088;
      20'h0a566: out <= 12'h088;
      20'h0a567: out <= 12'h088;
      20'h0a568: out <= 12'h088;
      20'h0a569: out <= 12'h088;
      20'h0a56a: out <= 12'h088;
      20'h0a56b: out <= 12'h088;
      20'h0a56c: out <= 12'h088;
      20'h0a56d: out <= 12'h088;
      20'h0a56e: out <= 12'h088;
      20'h0a56f: out <= 12'h088;
      20'h0a570: out <= 12'h088;
      20'h0a571: out <= 12'h088;
      20'h0a572: out <= 12'h088;
      20'h0a573: out <= 12'h088;
      20'h0a574: out <= 12'h088;
      20'h0a575: out <= 12'h088;
      20'h0a576: out <= 12'h088;
      20'h0a577: out <= 12'h088;
      20'h0a578: out <= 12'h088;
      20'h0a579: out <= 12'h088;
      20'h0a57a: out <= 12'h088;
      20'h0a57b: out <= 12'h088;
      20'h0a57c: out <= 12'h088;
      20'h0a57d: out <= 12'h088;
      20'h0a57e: out <= 12'h088;
      20'h0a57f: out <= 12'h088;
      20'h0a580: out <= 12'h088;
      20'h0a581: out <= 12'h088;
      20'h0a582: out <= 12'h088;
      20'h0a583: out <= 12'h088;
      20'h0a584: out <= 12'h088;
      20'h0a585: out <= 12'h088;
      20'h0a586: out <= 12'h088;
      20'h0a587: out <= 12'h088;
      20'h0a588: out <= 12'h088;
      20'h0a589: out <= 12'h088;
      20'h0a58a: out <= 12'h088;
      20'h0a58b: out <= 12'h088;
      20'h0a58c: out <= 12'h088;
      20'h0a58d: out <= 12'h088;
      20'h0a58e: out <= 12'h088;
      20'h0a58f: out <= 12'h088;
      20'h0a590: out <= 12'h088;
      20'h0a591: out <= 12'hee9;
      20'h0a592: out <= 12'hbb0;
      20'h0a593: out <= 12'h660;
      20'h0a594: out <= 12'h660;
      20'h0a595: out <= 12'h660;
      20'h0a596: out <= 12'h660;
      20'h0a597: out <= 12'h660;
      20'h0a598: out <= 12'h222;
      20'h0a599: out <= 12'h660;
      20'h0a59a: out <= 12'h660;
      20'h0a59b: out <= 12'h660;
      20'h0a59c: out <= 12'hee9;
      20'h0a59d: out <= 12'h660;
      20'h0a59e: out <= 12'hbb0;
      20'h0a59f: out <= 12'h660;
      20'h0a5a0: out <= 12'hbb0;
      20'h0a5a1: out <= 12'hee9;
      20'h0a5a2: out <= 12'hbb0;
      20'h0a5a3: out <= 12'h660;
      20'h0a5a4: out <= 12'h660;
      20'h0a5a5: out <= 12'h660;
      20'h0a5a6: out <= 12'hee9;
      20'h0a5a7: out <= 12'h660;
      20'h0a5a8: out <= 12'h603;
      20'h0a5a9: out <= 12'h603;
      20'h0a5aa: out <= 12'h603;
      20'h0a5ab: out <= 12'h603;
      20'h0a5ac: out <= 12'h000;
      20'h0a5ad: out <= 12'h000;
      20'h0a5ae: out <= 12'h000;
      20'h0a5af: out <= 12'h000;
      20'h0a5b0: out <= 12'h000;
      20'h0a5b1: out <= 12'h000;
      20'h0a5b2: out <= 12'h000;
      20'h0a5b3: out <= 12'h000;
      20'h0a5b4: out <= 12'h000;
      20'h0a5b5: out <= 12'h000;
      20'h0a5b6: out <= 12'h000;
      20'h0a5b7: out <= 12'h000;
      20'h0a5b8: out <= 12'h000;
      20'h0a5b9: out <= 12'h000;
      20'h0a5ba: out <= 12'h000;
      20'h0a5bb: out <= 12'h000;
      20'h0a5bc: out <= 12'h000;
      20'h0a5bd: out <= 12'h000;
      20'h0a5be: out <= 12'h000;
      20'h0a5bf: out <= 12'h000;
      20'h0a5c0: out <= 12'h000;
      20'h0a5c1: out <= 12'h000;
      20'h0a5c2: out <= 12'h000;
      20'h0a5c3: out <= 12'h000;
      20'h0a5c4: out <= 12'h000;
      20'h0a5c5: out <= 12'h000;
      20'h0a5c6: out <= 12'h000;
      20'h0a5c7: out <= 12'h000;
      20'h0a5c8: out <= 12'h000;
      20'h0a5c9: out <= 12'h000;
      20'h0a5ca: out <= 12'h000;
      20'h0a5cb: out <= 12'h000;
      20'h0a5cc: out <= 12'h000;
      20'h0a5cd: out <= 12'h000;
      20'h0a5ce: out <= 12'h000;
      20'h0a5cf: out <= 12'h000;
      20'h0a5d0: out <= 12'h000;
      20'h0a5d1: out <= 12'h000;
      20'h0a5d2: out <= 12'h000;
      20'h0a5d3: out <= 12'h000;
      20'h0a5d4: out <= 12'h000;
      20'h0a5d5: out <= 12'h000;
      20'h0a5d6: out <= 12'h000;
      20'h0a5d7: out <= 12'h000;
      20'h0a5d8: out <= 12'h000;
      20'h0a5d9: out <= 12'h000;
      20'h0a5da: out <= 12'h000;
      20'h0a5db: out <= 12'h000;
      20'h0a5dc: out <= 12'h000;
      20'h0a5dd: out <= 12'h000;
      20'h0a5de: out <= 12'h000;
      20'h0a5df: out <= 12'h000;
      20'h0a5e0: out <= 12'h000;
      20'h0a5e1: out <= 12'h000;
      20'h0a5e2: out <= 12'h000;
      20'h0a5e3: out <= 12'h000;
      20'h0a5e4: out <= 12'h000;
      20'h0a5e5: out <= 12'h000;
      20'h0a5e6: out <= 12'h000;
      20'h0a5e7: out <= 12'h000;
      20'h0a5e8: out <= 12'h000;
      20'h0a5e9: out <= 12'h000;
      20'h0a5ea: out <= 12'h000;
      20'h0a5eb: out <= 12'h000;
      20'h0a5ec: out <= 12'h000;
      20'h0a5ed: out <= 12'h000;
      20'h0a5ee: out <= 12'h000;
      20'h0a5ef: out <= 12'h000;
      20'h0a5f0: out <= 12'h000;
      20'h0a5f1: out <= 12'h000;
      20'h0a5f2: out <= 12'h000;
      20'h0a5f3: out <= 12'h000;
      20'h0a5f4: out <= 12'h000;
      20'h0a5f5: out <= 12'h000;
      20'h0a5f6: out <= 12'h000;
      20'h0a5f7: out <= 12'h000;
      20'h0a5f8: out <= 12'h000;
      20'h0a5f9: out <= 12'h000;
      20'h0a5fa: out <= 12'h000;
      20'h0a5fb: out <= 12'h000;
      20'h0a5fc: out <= 12'h603;
      20'h0a5fd: out <= 12'h603;
      20'h0a5fe: out <= 12'h603;
      20'h0a5ff: out <= 12'h603;
      20'h0a600: out <= 12'hb27;
      20'h0a601: out <= 12'hb27;
      20'h0a602: out <= 12'hb27;
      20'h0a603: out <= 12'hb27;
      20'h0a604: out <= 12'hb27;
      20'h0a605: out <= 12'hb27;
      20'h0a606: out <= 12'hb27;
      20'h0a607: out <= 12'hb27;
      20'h0a608: out <= 12'h000;
      20'h0a609: out <= 12'h000;
      20'h0a60a: out <= 12'h000;
      20'h0a60b: out <= 12'h000;
      20'h0a60c: out <= 12'h000;
      20'h0a60d: out <= 12'h000;
      20'h0a60e: out <= 12'h000;
      20'h0a60f: out <= 12'h000;
      20'h0a610: out <= 12'h000;
      20'h0a611: out <= 12'h000;
      20'h0a612: out <= 12'h000;
      20'h0a613: out <= 12'h000;
      20'h0a614: out <= 12'h000;
      20'h0a615: out <= 12'h000;
      20'h0a616: out <= 12'h000;
      20'h0a617: out <= 12'h000;
      20'h0a618: out <= 12'h000;
      20'h0a619: out <= 12'h000;
      20'h0a61a: out <= 12'h000;
      20'h0a61b: out <= 12'h000;
      20'h0a61c: out <= 12'h000;
      20'h0a61d: out <= 12'h000;
      20'h0a61e: out <= 12'h000;
      20'h0a61f: out <= 12'h000;
      20'h0a620: out <= 12'h000;
      20'h0a621: out <= 12'h000;
      20'h0a622: out <= 12'h000;
      20'h0a623: out <= 12'h000;
      20'h0a624: out <= 12'h000;
      20'h0a625: out <= 12'h000;
      20'h0a626: out <= 12'h000;
      20'h0a627: out <= 12'h000;
      20'h0a628: out <= 12'h4cd;
      20'h0a629: out <= 12'h4cd;
      20'h0a62a: out <= 12'h4cd;
      20'h0a62b: out <= 12'h4cd;
      20'h0a62c: out <= 12'h4cd;
      20'h0a62d: out <= 12'h4cd;
      20'h0a62e: out <= 12'h4cd;
      20'h0a62f: out <= 12'h4cd;
      20'h0a630: out <= 12'h5ef;
      20'h0a631: out <= 12'h5ef;
      20'h0a632: out <= 12'h5ef;
      20'h0a633: out <= 12'h5ef;
      20'h0a634: out <= 12'h5ef;
      20'h0a635: out <= 12'h5ef;
      20'h0a636: out <= 12'h5ef;
      20'h0a637: out <= 12'h5ef;
      20'h0a638: out <= 12'h000;
      20'h0a639: out <= 12'h000;
      20'h0a63a: out <= 12'h000;
      20'h0a63b: out <= 12'h000;
      20'h0a63c: out <= 12'h000;
      20'h0a63d: out <= 12'h000;
      20'h0a63e: out <= 12'h000;
      20'h0a63f: out <= 12'h000;
      20'h0a640: out <= 12'h088;
      20'h0a641: out <= 12'h088;
      20'h0a642: out <= 12'h088;
      20'h0a643: out <= 12'h088;
      20'h0a644: out <= 12'h088;
      20'h0a645: out <= 12'h088;
      20'h0a646: out <= 12'h088;
      20'h0a647: out <= 12'h088;
      20'h0a648: out <= 12'h088;
      20'h0a649: out <= 12'h088;
      20'h0a64a: out <= 12'h088;
      20'h0a64b: out <= 12'h088;
      20'h0a64c: out <= 12'h088;
      20'h0a64d: out <= 12'h088;
      20'h0a64e: out <= 12'h088;
      20'h0a64f: out <= 12'h088;
      20'h0a650: out <= 12'h088;
      20'h0a651: out <= 12'h088;
      20'h0a652: out <= 12'h088;
      20'h0a653: out <= 12'h088;
      20'h0a654: out <= 12'h088;
      20'h0a655: out <= 12'h088;
      20'h0a656: out <= 12'h088;
      20'h0a657: out <= 12'h088;
      20'h0a658: out <= 12'h088;
      20'h0a659: out <= 12'h088;
      20'h0a65a: out <= 12'h088;
      20'h0a65b: out <= 12'h088;
      20'h0a65c: out <= 12'h088;
      20'h0a65d: out <= 12'h088;
      20'h0a65e: out <= 12'h088;
      20'h0a65f: out <= 12'h088;
      20'h0a660: out <= 12'h088;
      20'h0a661: out <= 12'h088;
      20'h0a662: out <= 12'h088;
      20'h0a663: out <= 12'h088;
      20'h0a664: out <= 12'h088;
      20'h0a665: out <= 12'h088;
      20'h0a666: out <= 12'h088;
      20'h0a667: out <= 12'h088;
      20'h0a668: out <= 12'h088;
      20'h0a669: out <= 12'h088;
      20'h0a66a: out <= 12'h088;
      20'h0a66b: out <= 12'h088;
      20'h0a66c: out <= 12'h088;
      20'h0a66d: out <= 12'h088;
      20'h0a66e: out <= 12'h088;
      20'h0a66f: out <= 12'h088;
      20'h0a670: out <= 12'h088;
      20'h0a671: out <= 12'h088;
      20'h0a672: out <= 12'h088;
      20'h0a673: out <= 12'h088;
      20'h0a674: out <= 12'h088;
      20'h0a675: out <= 12'h088;
      20'h0a676: out <= 12'h088;
      20'h0a677: out <= 12'h088;
      20'h0a678: out <= 12'h088;
      20'h0a679: out <= 12'h088;
      20'h0a67a: out <= 12'h088;
      20'h0a67b: out <= 12'h088;
      20'h0a67c: out <= 12'h088;
      20'h0a67d: out <= 12'h088;
      20'h0a67e: out <= 12'h088;
      20'h0a67f: out <= 12'h088;
      20'h0a680: out <= 12'h088;
      20'h0a681: out <= 12'h088;
      20'h0a682: out <= 12'h088;
      20'h0a683: out <= 12'h088;
      20'h0a684: out <= 12'h088;
      20'h0a685: out <= 12'h088;
      20'h0a686: out <= 12'h088;
      20'h0a687: out <= 12'h088;
      20'h0a688: out <= 12'h088;
      20'h0a689: out <= 12'h088;
      20'h0a68a: out <= 12'h088;
      20'h0a68b: out <= 12'h088;
      20'h0a68c: out <= 12'h088;
      20'h0a68d: out <= 12'h088;
      20'h0a68e: out <= 12'h088;
      20'h0a68f: out <= 12'h088;
      20'h0a690: out <= 12'h088;
      20'h0a691: out <= 12'h088;
      20'h0a692: out <= 12'h088;
      20'h0a693: out <= 12'h088;
      20'h0a694: out <= 12'h088;
      20'h0a695: out <= 12'h088;
      20'h0a696: out <= 12'h088;
      20'h0a697: out <= 12'h088;
      20'h0a698: out <= 12'h088;
      20'h0a699: out <= 12'h088;
      20'h0a69a: out <= 12'h088;
      20'h0a69b: out <= 12'h088;
      20'h0a69c: out <= 12'h088;
      20'h0a69d: out <= 12'h088;
      20'h0a69e: out <= 12'h088;
      20'h0a69f: out <= 12'h088;
      20'h0a6a0: out <= 12'h088;
      20'h0a6a1: out <= 12'h088;
      20'h0a6a2: out <= 12'h088;
      20'h0a6a3: out <= 12'h088;
      20'h0a6a4: out <= 12'h088;
      20'h0a6a5: out <= 12'h088;
      20'h0a6a6: out <= 12'h088;
      20'h0a6a7: out <= 12'h088;
      20'h0a6a8: out <= 12'h088;
      20'h0a6a9: out <= 12'h660;
      20'h0a6aa: out <= 12'hbb0;
      20'h0a6ab: out <= 12'h660;
      20'h0a6ac: out <= 12'h660;
      20'h0a6ad: out <= 12'h660;
      20'h0a6ae: out <= 12'hee9;
      20'h0a6af: out <= 12'h660;
      20'h0a6b0: out <= 12'h222;
      20'h0a6b1: out <= 12'h660;
      20'h0a6b2: out <= 12'hee9;
      20'h0a6b3: out <= 12'h660;
      20'h0a6b4: out <= 12'hee9;
      20'h0a6b5: out <= 12'h660;
      20'h0a6b6: out <= 12'hbb0;
      20'h0a6b7: out <= 12'h660;
      20'h0a6b8: out <= 12'h660;
      20'h0a6b9: out <= 12'h660;
      20'h0a6ba: out <= 12'hbb0;
      20'h0a6bb: out <= 12'h660;
      20'h0a6bc: out <= 12'h660;
      20'h0a6bd: out <= 12'h660;
      20'h0a6be: out <= 12'h660;
      20'h0a6bf: out <= 12'h660;
      20'h0a6c0: out <= 12'h603;
      20'h0a6c1: out <= 12'h603;
      20'h0a6c2: out <= 12'h603;
      20'h0a6c3: out <= 12'h603;
      20'h0a6c4: out <= 12'h000;
      20'h0a6c5: out <= 12'hbbb;
      20'h0a6c6: out <= 12'hbbb;
      20'h0a6c7: out <= 12'hbbb;
      20'h0a6c8: out <= 12'hbbb;
      20'h0a6c9: out <= 12'hbbb;
      20'h0a6ca: out <= 12'h000;
      20'h0a6cb: out <= 12'h000;
      20'h0a6cc: out <= 12'h000;
      20'h0a6cd: out <= 12'h000;
      20'h0a6ce: out <= 12'h000;
      20'h0a6cf: out <= 12'hbbb;
      20'h0a6d0: out <= 12'hbbb;
      20'h0a6d1: out <= 12'h000;
      20'h0a6d2: out <= 12'h000;
      20'h0a6d3: out <= 12'h000;
      20'h0a6d4: out <= 12'h000;
      20'h0a6d5: out <= 12'hbbb;
      20'h0a6d6: out <= 12'hbbb;
      20'h0a6d7: out <= 12'hbbb;
      20'h0a6d8: out <= 12'hbbb;
      20'h0a6d9: out <= 12'hbbb;
      20'h0a6da: out <= 12'h000;
      20'h0a6db: out <= 12'h000;
      20'h0a6dc: out <= 12'h000;
      20'h0a6dd: out <= 12'hbbb;
      20'h0a6de: out <= 12'hbbb;
      20'h0a6df: out <= 12'hbbb;
      20'h0a6e0: out <= 12'hbbb;
      20'h0a6e1: out <= 12'hbbb;
      20'h0a6e2: out <= 12'h000;
      20'h0a6e3: out <= 12'h000;
      20'h0a6e4: out <= 12'h000;
      20'h0a6e5: out <= 12'h000;
      20'h0a6e6: out <= 12'h000;
      20'h0a6e7: out <= 12'hbbb;
      20'h0a6e8: out <= 12'hbbb;
      20'h0a6e9: out <= 12'hbbb;
      20'h0a6ea: out <= 12'h000;
      20'h0a6eb: out <= 12'h000;
      20'h0a6ec: out <= 12'hbbb;
      20'h0a6ed: out <= 12'hbbb;
      20'h0a6ee: out <= 12'hbbb;
      20'h0a6ef: out <= 12'hbbb;
      20'h0a6f0: out <= 12'hbbb;
      20'h0a6f1: out <= 12'hbbb;
      20'h0a6f2: out <= 12'hbbb;
      20'h0a6f3: out <= 12'h000;
      20'h0a6f4: out <= 12'h000;
      20'h0a6f5: out <= 12'h000;
      20'h0a6f6: out <= 12'hbbb;
      20'h0a6f7: out <= 12'hbbb;
      20'h0a6f8: out <= 12'hbbb;
      20'h0a6f9: out <= 12'hbbb;
      20'h0a6fa: out <= 12'h000;
      20'h0a6fb: out <= 12'h000;
      20'h0a6fc: out <= 12'hbbb;
      20'h0a6fd: out <= 12'hbbb;
      20'h0a6fe: out <= 12'hbbb;
      20'h0a6ff: out <= 12'hbbb;
      20'h0a700: out <= 12'hbbb;
      20'h0a701: out <= 12'hbbb;
      20'h0a702: out <= 12'hbbb;
      20'h0a703: out <= 12'h000;
      20'h0a704: out <= 12'h000;
      20'h0a705: out <= 12'hbbb;
      20'h0a706: out <= 12'hbbb;
      20'h0a707: out <= 12'hbbb;
      20'h0a708: out <= 12'hbbb;
      20'h0a709: out <= 12'hbbb;
      20'h0a70a: out <= 12'h000;
      20'h0a70b: out <= 12'h000;
      20'h0a70c: out <= 12'h000;
      20'h0a70d: out <= 12'hbbb;
      20'h0a70e: out <= 12'hbbb;
      20'h0a70f: out <= 12'hbbb;
      20'h0a710: out <= 12'hbbb;
      20'h0a711: out <= 12'hbbb;
      20'h0a712: out <= 12'h000;
      20'h0a713: out <= 12'h000;
      20'h0a714: out <= 12'h603;
      20'h0a715: out <= 12'h603;
      20'h0a716: out <= 12'h603;
      20'h0a717: out <= 12'h603;
      20'h0a718: out <= 12'hee9;
      20'h0a719: out <= 12'hee9;
      20'h0a71a: out <= 12'hee9;
      20'h0a71b: out <= 12'hee9;
      20'h0a71c: out <= 12'hee9;
      20'h0a71d: out <= 12'hee9;
      20'h0a71e: out <= 12'hee9;
      20'h0a71f: out <= 12'hb27;
      20'h0a720: out <= 12'h000;
      20'h0a721: out <= 12'h000;
      20'h0a722: out <= 12'h000;
      20'h0a723: out <= 12'h000;
      20'h0a724: out <= 12'h000;
      20'h0a725: out <= 12'h000;
      20'h0a726: out <= 12'h000;
      20'h0a727: out <= 12'h000;
      20'h0a728: out <= 12'hfa9;
      20'h0a729: out <= 12'hfa9;
      20'h0a72a: out <= 12'hfa9;
      20'h0a72b: out <= 12'hfa9;
      20'h0a72c: out <= 12'hfa9;
      20'h0a72d: out <= 12'hfa9;
      20'h0a72e: out <= 12'hfa9;
      20'h0a72f: out <= 12'hfa9;
      20'h0a730: out <= 12'hf76;
      20'h0a731: out <= 12'hf76;
      20'h0a732: out <= 12'hf76;
      20'h0a733: out <= 12'hf76;
      20'h0a734: out <= 12'hf76;
      20'h0a735: out <= 12'hf76;
      20'h0a736: out <= 12'hf76;
      20'h0a737: out <= 12'hf76;
      20'h0a738: out <= 12'hfa9;
      20'h0a739: out <= 12'hfa9;
      20'h0a73a: out <= 12'hfa9;
      20'h0a73b: out <= 12'hfa9;
      20'h0a73c: out <= 12'hfa9;
      20'h0a73d: out <= 12'hfa9;
      20'h0a73e: out <= 12'hfa9;
      20'h0a73f: out <= 12'hfa9;
      20'h0a740: out <= 12'hf76;
      20'h0a741: out <= 12'hf76;
      20'h0a742: out <= 12'hf76;
      20'h0a743: out <= 12'hf76;
      20'h0a744: out <= 12'hf76;
      20'h0a745: out <= 12'hf76;
      20'h0a746: out <= 12'hf76;
      20'h0a747: out <= 12'hf76;
      20'h0a748: out <= 12'hfa9;
      20'h0a749: out <= 12'hfa9;
      20'h0a74a: out <= 12'hfa9;
      20'h0a74b: out <= 12'hfa9;
      20'h0a74c: out <= 12'hfa9;
      20'h0a74d: out <= 12'hfa9;
      20'h0a74e: out <= 12'hfa9;
      20'h0a74f: out <= 12'hfa9;
      20'h0a750: out <= 12'h000;
      20'h0a751: out <= 12'h000;
      20'h0a752: out <= 12'h000;
      20'h0a753: out <= 12'h000;
      20'h0a754: out <= 12'h000;
      20'h0a755: out <= 12'h000;
      20'h0a756: out <= 12'h000;
      20'h0a757: out <= 12'h000;
      20'h0a758: out <= 12'h088;
      20'h0a759: out <= 12'h088;
      20'h0a75a: out <= 12'h088;
      20'h0a75b: out <= 12'h088;
      20'h0a75c: out <= 12'h088;
      20'h0a75d: out <= 12'h088;
      20'h0a75e: out <= 12'h088;
      20'h0a75f: out <= 12'h088;
      20'h0a760: out <= 12'h088;
      20'h0a761: out <= 12'h088;
      20'h0a762: out <= 12'h088;
      20'h0a763: out <= 12'h088;
      20'h0a764: out <= 12'h088;
      20'h0a765: out <= 12'h088;
      20'h0a766: out <= 12'h088;
      20'h0a767: out <= 12'h088;
      20'h0a768: out <= 12'h088;
      20'h0a769: out <= 12'h088;
      20'h0a76a: out <= 12'h088;
      20'h0a76b: out <= 12'h088;
      20'h0a76c: out <= 12'h088;
      20'h0a76d: out <= 12'h088;
      20'h0a76e: out <= 12'h088;
      20'h0a76f: out <= 12'h088;
      20'h0a770: out <= 12'h088;
      20'h0a771: out <= 12'h088;
      20'h0a772: out <= 12'h088;
      20'h0a773: out <= 12'h088;
      20'h0a774: out <= 12'h088;
      20'h0a775: out <= 12'h088;
      20'h0a776: out <= 12'h088;
      20'h0a777: out <= 12'h088;
      20'h0a778: out <= 12'h088;
      20'h0a779: out <= 12'h088;
      20'h0a77a: out <= 12'h088;
      20'h0a77b: out <= 12'h088;
      20'h0a77c: out <= 12'h088;
      20'h0a77d: out <= 12'h088;
      20'h0a77e: out <= 12'h088;
      20'h0a77f: out <= 12'h088;
      20'h0a780: out <= 12'h088;
      20'h0a781: out <= 12'h088;
      20'h0a782: out <= 12'h088;
      20'h0a783: out <= 12'h088;
      20'h0a784: out <= 12'h088;
      20'h0a785: out <= 12'h088;
      20'h0a786: out <= 12'h088;
      20'h0a787: out <= 12'h088;
      20'h0a788: out <= 12'h088;
      20'h0a789: out <= 12'h088;
      20'h0a78a: out <= 12'h088;
      20'h0a78b: out <= 12'h088;
      20'h0a78c: out <= 12'h088;
      20'h0a78d: out <= 12'h088;
      20'h0a78e: out <= 12'h088;
      20'h0a78f: out <= 12'h088;
      20'h0a790: out <= 12'h088;
      20'h0a791: out <= 12'h088;
      20'h0a792: out <= 12'h088;
      20'h0a793: out <= 12'h088;
      20'h0a794: out <= 12'h088;
      20'h0a795: out <= 12'h088;
      20'h0a796: out <= 12'h088;
      20'h0a797: out <= 12'h088;
      20'h0a798: out <= 12'h088;
      20'h0a799: out <= 12'h088;
      20'h0a79a: out <= 12'h088;
      20'h0a79b: out <= 12'h088;
      20'h0a79c: out <= 12'h088;
      20'h0a79d: out <= 12'h088;
      20'h0a79e: out <= 12'h088;
      20'h0a79f: out <= 12'h088;
      20'h0a7a0: out <= 12'h088;
      20'h0a7a1: out <= 12'h088;
      20'h0a7a2: out <= 12'h088;
      20'h0a7a3: out <= 12'h088;
      20'h0a7a4: out <= 12'h088;
      20'h0a7a5: out <= 12'h088;
      20'h0a7a6: out <= 12'h088;
      20'h0a7a7: out <= 12'h088;
      20'h0a7a8: out <= 12'h088;
      20'h0a7a9: out <= 12'h088;
      20'h0a7aa: out <= 12'h088;
      20'h0a7ab: out <= 12'h088;
      20'h0a7ac: out <= 12'h088;
      20'h0a7ad: out <= 12'h088;
      20'h0a7ae: out <= 12'h088;
      20'h0a7af: out <= 12'h088;
      20'h0a7b0: out <= 12'h088;
      20'h0a7b1: out <= 12'h088;
      20'h0a7b2: out <= 12'h088;
      20'h0a7b3: out <= 12'h088;
      20'h0a7b4: out <= 12'h088;
      20'h0a7b5: out <= 12'h088;
      20'h0a7b6: out <= 12'h088;
      20'h0a7b7: out <= 12'h088;
      20'h0a7b8: out <= 12'h088;
      20'h0a7b9: out <= 12'h088;
      20'h0a7ba: out <= 12'h088;
      20'h0a7bb: out <= 12'h088;
      20'h0a7bc: out <= 12'h088;
      20'h0a7bd: out <= 12'h088;
      20'h0a7be: out <= 12'h088;
      20'h0a7bf: out <= 12'h088;
      20'h0a7c0: out <= 12'h088;
      20'h0a7c1: out <= 12'hbb0;
      20'h0a7c2: out <= 12'hbb0;
      20'h0a7c3: out <= 12'h660;
      20'h0a7c4: out <= 12'h660;
      20'h0a7c5: out <= 12'h660;
      20'h0a7c6: out <= 12'h660;
      20'h0a7c7: out <= 12'h660;
      20'h0a7c8: out <= 12'h222;
      20'h0a7c9: out <= 12'h660;
      20'h0a7ca: out <= 12'h660;
      20'h0a7cb: out <= 12'h660;
      20'h0a7cc: out <= 12'hee9;
      20'h0a7cd: out <= 12'h660;
      20'h0a7ce: out <= 12'hbb0;
      20'h0a7cf: out <= 12'hbb0;
      20'h0a7d0: out <= 12'hbb0;
      20'h0a7d1: out <= 12'hbb0;
      20'h0a7d2: out <= 12'hbb0;
      20'h0a7d3: out <= 12'h660;
      20'h0a7d4: out <= 12'h660;
      20'h0a7d5: out <= 12'h660;
      20'h0a7d6: out <= 12'hee9;
      20'h0a7d7: out <= 12'h660;
      20'h0a7d8: out <= 12'h603;
      20'h0a7d9: out <= 12'h603;
      20'h0a7da: out <= 12'h603;
      20'h0a7db: out <= 12'h603;
      20'h0a7dc: out <= 12'hbbb;
      20'h0a7dd: out <= 12'hbbb;
      20'h0a7de: out <= 12'h000;
      20'h0a7df: out <= 12'h000;
      20'h0a7e0: out <= 12'h000;
      20'h0a7e1: out <= 12'hbbb;
      20'h0a7e2: out <= 12'hbbb;
      20'h0a7e3: out <= 12'h000;
      20'h0a7e4: out <= 12'h000;
      20'h0a7e5: out <= 12'h000;
      20'h0a7e6: out <= 12'hbbb;
      20'h0a7e7: out <= 12'hbbb;
      20'h0a7e8: out <= 12'hbbb;
      20'h0a7e9: out <= 12'h000;
      20'h0a7ea: out <= 12'h000;
      20'h0a7eb: out <= 12'h000;
      20'h0a7ec: out <= 12'hbbb;
      20'h0a7ed: out <= 12'hbbb;
      20'h0a7ee: out <= 12'h000;
      20'h0a7ef: out <= 12'h000;
      20'h0a7f0: out <= 12'h000;
      20'h0a7f1: out <= 12'hbbb;
      20'h0a7f2: out <= 12'hbbb;
      20'h0a7f3: out <= 12'h000;
      20'h0a7f4: out <= 12'hbbb;
      20'h0a7f5: out <= 12'hbbb;
      20'h0a7f6: out <= 12'h000;
      20'h0a7f7: out <= 12'h000;
      20'h0a7f8: out <= 12'h000;
      20'h0a7f9: out <= 12'hbbb;
      20'h0a7fa: out <= 12'hbbb;
      20'h0a7fb: out <= 12'h000;
      20'h0a7fc: out <= 12'h000;
      20'h0a7fd: out <= 12'h000;
      20'h0a7fe: out <= 12'hbbb;
      20'h0a7ff: out <= 12'hbbb;
      20'h0a800: out <= 12'hbbb;
      20'h0a801: out <= 12'hbbb;
      20'h0a802: out <= 12'h000;
      20'h0a803: out <= 12'h000;
      20'h0a804: out <= 12'hbbb;
      20'h0a805: out <= 12'hbbb;
      20'h0a806: out <= 12'h000;
      20'h0a807: out <= 12'h000;
      20'h0a808: out <= 12'h000;
      20'h0a809: out <= 12'h000;
      20'h0a80a: out <= 12'h000;
      20'h0a80b: out <= 12'h000;
      20'h0a80c: out <= 12'h000;
      20'h0a80d: out <= 12'hbbb;
      20'h0a80e: out <= 12'hbbb;
      20'h0a80f: out <= 12'h000;
      20'h0a810: out <= 12'h000;
      20'h0a811: out <= 12'h000;
      20'h0a812: out <= 12'h000;
      20'h0a813: out <= 12'h000;
      20'h0a814: out <= 12'hbbb;
      20'h0a815: out <= 12'hbbb;
      20'h0a816: out <= 12'h000;
      20'h0a817: out <= 12'h000;
      20'h0a818: out <= 12'h000;
      20'h0a819: out <= 12'hbbb;
      20'h0a81a: out <= 12'hbbb;
      20'h0a81b: out <= 12'h000;
      20'h0a81c: out <= 12'hbbb;
      20'h0a81d: out <= 12'hbbb;
      20'h0a81e: out <= 12'h000;
      20'h0a81f: out <= 12'h000;
      20'h0a820: out <= 12'h000;
      20'h0a821: out <= 12'hbbb;
      20'h0a822: out <= 12'hbbb;
      20'h0a823: out <= 12'h000;
      20'h0a824: out <= 12'hbbb;
      20'h0a825: out <= 12'hbbb;
      20'h0a826: out <= 12'h000;
      20'h0a827: out <= 12'h000;
      20'h0a828: out <= 12'h000;
      20'h0a829: out <= 12'hbbb;
      20'h0a82a: out <= 12'hbbb;
      20'h0a82b: out <= 12'h000;
      20'h0a82c: out <= 12'h603;
      20'h0a82d: out <= 12'h603;
      20'h0a82e: out <= 12'h603;
      20'h0a82f: out <= 12'h603;
      20'h0a830: out <= 12'hee9;
      20'h0a831: out <= 12'hf87;
      20'h0a832: out <= 12'hf87;
      20'h0a833: out <= 12'hf87;
      20'h0a834: out <= 12'hf87;
      20'h0a835: out <= 12'hf87;
      20'h0a836: out <= 12'hf87;
      20'h0a837: out <= 12'hb27;
      20'h0a838: out <= 12'h000;
      20'h0a839: out <= 12'h000;
      20'h0a83a: out <= 12'h000;
      20'h0a83b: out <= 12'h000;
      20'h0a83c: out <= 12'h000;
      20'h0a83d: out <= 12'h000;
      20'h0a83e: out <= 12'h000;
      20'h0a83f: out <= 12'h000;
      20'h0a840: out <= 12'hfa9;
      20'h0a841: out <= 12'hfa9;
      20'h0a842: out <= 12'hfa9;
      20'h0a843: out <= 12'hfa9;
      20'h0a844: out <= 12'hfa9;
      20'h0a845: out <= 12'hfa9;
      20'h0a846: out <= 12'hfa9;
      20'h0a847: out <= 12'hfa9;
      20'h0a848: out <= 12'hf76;
      20'h0a849: out <= 12'hf76;
      20'h0a84a: out <= 12'hf76;
      20'h0a84b: out <= 12'hf76;
      20'h0a84c: out <= 12'hf76;
      20'h0a84d: out <= 12'hf76;
      20'h0a84e: out <= 12'hf76;
      20'h0a84f: out <= 12'hf76;
      20'h0a850: out <= 12'hfa9;
      20'h0a851: out <= 12'hfa9;
      20'h0a852: out <= 12'hfa9;
      20'h0a853: out <= 12'hfa9;
      20'h0a854: out <= 12'hfa9;
      20'h0a855: out <= 12'hfa9;
      20'h0a856: out <= 12'hfa9;
      20'h0a857: out <= 12'hfa9;
      20'h0a858: out <= 12'hf76;
      20'h0a859: out <= 12'hf76;
      20'h0a85a: out <= 12'hf76;
      20'h0a85b: out <= 12'hf76;
      20'h0a85c: out <= 12'hf76;
      20'h0a85d: out <= 12'hf76;
      20'h0a85e: out <= 12'hf76;
      20'h0a85f: out <= 12'hf76;
      20'h0a860: out <= 12'hfa9;
      20'h0a861: out <= 12'hfa9;
      20'h0a862: out <= 12'hfa9;
      20'h0a863: out <= 12'hfa9;
      20'h0a864: out <= 12'hfa9;
      20'h0a865: out <= 12'hfa9;
      20'h0a866: out <= 12'hfa9;
      20'h0a867: out <= 12'hfa9;
      20'h0a868: out <= 12'h000;
      20'h0a869: out <= 12'h000;
      20'h0a86a: out <= 12'h000;
      20'h0a86b: out <= 12'h000;
      20'h0a86c: out <= 12'h000;
      20'h0a86d: out <= 12'h000;
      20'h0a86e: out <= 12'h000;
      20'h0a86f: out <= 12'h000;
      20'h0a870: out <= 12'h088;
      20'h0a871: out <= 12'h088;
      20'h0a872: out <= 12'h088;
      20'h0a873: out <= 12'h088;
      20'h0a874: out <= 12'h088;
      20'h0a875: out <= 12'h088;
      20'h0a876: out <= 12'h088;
      20'h0a877: out <= 12'h088;
      20'h0a878: out <= 12'h088;
      20'h0a879: out <= 12'h088;
      20'h0a87a: out <= 12'h088;
      20'h0a87b: out <= 12'h088;
      20'h0a87c: out <= 12'h088;
      20'h0a87d: out <= 12'h088;
      20'h0a87e: out <= 12'h088;
      20'h0a87f: out <= 12'h088;
      20'h0a880: out <= 12'h088;
      20'h0a881: out <= 12'h088;
      20'h0a882: out <= 12'h088;
      20'h0a883: out <= 12'h088;
      20'h0a884: out <= 12'h088;
      20'h0a885: out <= 12'h088;
      20'h0a886: out <= 12'h088;
      20'h0a887: out <= 12'h088;
      20'h0a888: out <= 12'h088;
      20'h0a889: out <= 12'h088;
      20'h0a88a: out <= 12'h088;
      20'h0a88b: out <= 12'h088;
      20'h0a88c: out <= 12'h088;
      20'h0a88d: out <= 12'h088;
      20'h0a88e: out <= 12'h088;
      20'h0a88f: out <= 12'h088;
      20'h0a890: out <= 12'h088;
      20'h0a891: out <= 12'h088;
      20'h0a892: out <= 12'h088;
      20'h0a893: out <= 12'h088;
      20'h0a894: out <= 12'h088;
      20'h0a895: out <= 12'h088;
      20'h0a896: out <= 12'h088;
      20'h0a897: out <= 12'h088;
      20'h0a898: out <= 12'h088;
      20'h0a899: out <= 12'h088;
      20'h0a89a: out <= 12'h088;
      20'h0a89b: out <= 12'h088;
      20'h0a89c: out <= 12'h088;
      20'h0a89d: out <= 12'h088;
      20'h0a89e: out <= 12'h088;
      20'h0a89f: out <= 12'h088;
      20'h0a8a0: out <= 12'h088;
      20'h0a8a1: out <= 12'h088;
      20'h0a8a2: out <= 12'h088;
      20'h0a8a3: out <= 12'h088;
      20'h0a8a4: out <= 12'h088;
      20'h0a8a5: out <= 12'h088;
      20'h0a8a6: out <= 12'h088;
      20'h0a8a7: out <= 12'h088;
      20'h0a8a8: out <= 12'h088;
      20'h0a8a9: out <= 12'h088;
      20'h0a8aa: out <= 12'h088;
      20'h0a8ab: out <= 12'h088;
      20'h0a8ac: out <= 12'h088;
      20'h0a8ad: out <= 12'h088;
      20'h0a8ae: out <= 12'h088;
      20'h0a8af: out <= 12'h088;
      20'h0a8b0: out <= 12'h088;
      20'h0a8b1: out <= 12'h088;
      20'h0a8b2: out <= 12'h088;
      20'h0a8b3: out <= 12'h088;
      20'h0a8b4: out <= 12'h088;
      20'h0a8b5: out <= 12'h088;
      20'h0a8b6: out <= 12'h088;
      20'h0a8b7: out <= 12'h088;
      20'h0a8b8: out <= 12'h088;
      20'h0a8b9: out <= 12'h088;
      20'h0a8ba: out <= 12'h088;
      20'h0a8bb: out <= 12'h088;
      20'h0a8bc: out <= 12'h088;
      20'h0a8bd: out <= 12'h088;
      20'h0a8be: out <= 12'h088;
      20'h0a8bf: out <= 12'h088;
      20'h0a8c0: out <= 12'h088;
      20'h0a8c1: out <= 12'h088;
      20'h0a8c2: out <= 12'h088;
      20'h0a8c3: out <= 12'h088;
      20'h0a8c4: out <= 12'h088;
      20'h0a8c5: out <= 12'h088;
      20'h0a8c6: out <= 12'h088;
      20'h0a8c7: out <= 12'h088;
      20'h0a8c8: out <= 12'h088;
      20'h0a8c9: out <= 12'h088;
      20'h0a8ca: out <= 12'h088;
      20'h0a8cb: out <= 12'h088;
      20'h0a8cc: out <= 12'h088;
      20'h0a8cd: out <= 12'h088;
      20'h0a8ce: out <= 12'h088;
      20'h0a8cf: out <= 12'h088;
      20'h0a8d0: out <= 12'h088;
      20'h0a8d1: out <= 12'h088;
      20'h0a8d2: out <= 12'h088;
      20'h0a8d3: out <= 12'h088;
      20'h0a8d4: out <= 12'h088;
      20'h0a8d5: out <= 12'h088;
      20'h0a8d6: out <= 12'h088;
      20'h0a8d7: out <= 12'h088;
      20'h0a8d8: out <= 12'h088;
      20'h0a8d9: out <= 12'h660;
      20'h0a8da: out <= 12'h660;
      20'h0a8db: out <= 12'h660;
      20'h0a8dc: out <= 12'h660;
      20'h0a8dd: out <= 12'h660;
      20'h0a8de: out <= 12'hee9;
      20'h0a8df: out <= 12'h660;
      20'h0a8e0: out <= 12'h222;
      20'h0a8e1: out <= 12'h660;
      20'h0a8e2: out <= 12'hee9;
      20'h0a8e3: out <= 12'h660;
      20'h0a8e4: out <= 12'hee9;
      20'h0a8e5: out <= 12'h660;
      20'h0a8e6: out <= 12'h660;
      20'h0a8e7: out <= 12'h660;
      20'h0a8e8: out <= 12'h660;
      20'h0a8e9: out <= 12'h660;
      20'h0a8ea: out <= 12'h660;
      20'h0a8eb: out <= 12'h660;
      20'h0a8ec: out <= 12'h660;
      20'h0a8ed: out <= 12'h660;
      20'h0a8ee: out <= 12'h660;
      20'h0a8ef: out <= 12'h660;
      20'h0a8f0: out <= 12'h603;
      20'h0a8f1: out <= 12'h603;
      20'h0a8f2: out <= 12'h603;
      20'h0a8f3: out <= 12'h603;
      20'h0a8f4: out <= 12'hbbb;
      20'h0a8f5: out <= 12'hbbb;
      20'h0a8f6: out <= 12'h000;
      20'h0a8f7: out <= 12'h000;
      20'h0a8f8: out <= 12'hbbb;
      20'h0a8f9: out <= 12'hbbb;
      20'h0a8fa: out <= 12'hbbb;
      20'h0a8fb: out <= 12'h000;
      20'h0a8fc: out <= 12'h000;
      20'h0a8fd: out <= 12'h000;
      20'h0a8fe: out <= 12'h000;
      20'h0a8ff: out <= 12'hbbb;
      20'h0a900: out <= 12'hbbb;
      20'h0a901: out <= 12'h000;
      20'h0a902: out <= 12'h000;
      20'h0a903: out <= 12'h000;
      20'h0a904: out <= 12'h000;
      20'h0a905: out <= 12'h000;
      20'h0a906: out <= 12'h000;
      20'h0a907: out <= 12'h000;
      20'h0a908: out <= 12'h000;
      20'h0a909: out <= 12'hbbb;
      20'h0a90a: out <= 12'hbbb;
      20'h0a90b: out <= 12'h000;
      20'h0a90c: out <= 12'h000;
      20'h0a90d: out <= 12'h000;
      20'h0a90e: out <= 12'h000;
      20'h0a90f: out <= 12'h000;
      20'h0a910: out <= 12'h000;
      20'h0a911: out <= 12'hbbb;
      20'h0a912: out <= 12'hbbb;
      20'h0a913: out <= 12'h000;
      20'h0a914: out <= 12'h000;
      20'h0a915: out <= 12'hbbb;
      20'h0a916: out <= 12'hbbb;
      20'h0a917: out <= 12'h000;
      20'h0a918: out <= 12'hbbb;
      20'h0a919: out <= 12'hbbb;
      20'h0a91a: out <= 12'h000;
      20'h0a91b: out <= 12'h000;
      20'h0a91c: out <= 12'hbbb;
      20'h0a91d: out <= 12'hbbb;
      20'h0a91e: out <= 12'hbbb;
      20'h0a91f: out <= 12'hbbb;
      20'h0a920: out <= 12'hbbb;
      20'h0a921: out <= 12'hbbb;
      20'h0a922: out <= 12'h000;
      20'h0a923: out <= 12'h000;
      20'h0a924: out <= 12'hbbb;
      20'h0a925: out <= 12'hbbb;
      20'h0a926: out <= 12'h000;
      20'h0a927: out <= 12'h000;
      20'h0a928: out <= 12'h000;
      20'h0a929: out <= 12'h000;
      20'h0a92a: out <= 12'h000;
      20'h0a92b: out <= 12'h000;
      20'h0a92c: out <= 12'h000;
      20'h0a92d: out <= 12'h000;
      20'h0a92e: out <= 12'h000;
      20'h0a92f: out <= 12'h000;
      20'h0a930: out <= 12'hbbb;
      20'h0a931: out <= 12'hbbb;
      20'h0a932: out <= 12'h000;
      20'h0a933: out <= 12'h000;
      20'h0a934: out <= 12'hbbb;
      20'h0a935: out <= 12'hbbb;
      20'h0a936: out <= 12'h000;
      20'h0a937: out <= 12'h000;
      20'h0a938: out <= 12'h000;
      20'h0a939: out <= 12'hbbb;
      20'h0a93a: out <= 12'hbbb;
      20'h0a93b: out <= 12'h000;
      20'h0a93c: out <= 12'hbbb;
      20'h0a93d: out <= 12'hbbb;
      20'h0a93e: out <= 12'h000;
      20'h0a93f: out <= 12'h000;
      20'h0a940: out <= 12'h000;
      20'h0a941: out <= 12'hbbb;
      20'h0a942: out <= 12'hbbb;
      20'h0a943: out <= 12'h000;
      20'h0a944: out <= 12'h603;
      20'h0a945: out <= 12'h603;
      20'h0a946: out <= 12'h603;
      20'h0a947: out <= 12'h603;
      20'h0a948: out <= 12'hee9;
      20'h0a949: out <= 12'hf87;
      20'h0a94a: out <= 12'hee9;
      20'h0a94b: out <= 12'hee9;
      20'h0a94c: out <= 12'hee9;
      20'h0a94d: out <= 12'hb27;
      20'h0a94e: out <= 12'hf87;
      20'h0a94f: out <= 12'hb27;
      20'h0a950: out <= 12'h000;
      20'h0a951: out <= 12'h000;
      20'h0a952: out <= 12'h000;
      20'h0a953: out <= 12'h000;
      20'h0a954: out <= 12'h000;
      20'h0a955: out <= 12'h000;
      20'h0a956: out <= 12'h000;
      20'h0a957: out <= 12'h000;
      20'h0a958: out <= 12'hfa9;
      20'h0a959: out <= 12'hfa9;
      20'h0a95a: out <= 12'hfa9;
      20'h0a95b: out <= 12'hfa9;
      20'h0a95c: out <= 12'hfa9;
      20'h0a95d: out <= 12'hfa9;
      20'h0a95e: out <= 12'hfa9;
      20'h0a95f: out <= 12'hfa9;
      20'h0a960: out <= 12'hf76;
      20'h0a961: out <= 12'hf76;
      20'h0a962: out <= 12'hf76;
      20'h0a963: out <= 12'hf76;
      20'h0a964: out <= 12'hf76;
      20'h0a965: out <= 12'hf76;
      20'h0a966: out <= 12'hf76;
      20'h0a967: out <= 12'hf76;
      20'h0a968: out <= 12'hfa9;
      20'h0a969: out <= 12'hfa9;
      20'h0a96a: out <= 12'hfa9;
      20'h0a96b: out <= 12'hfa9;
      20'h0a96c: out <= 12'hfa9;
      20'h0a96d: out <= 12'hfa9;
      20'h0a96e: out <= 12'hfa9;
      20'h0a96f: out <= 12'hfa9;
      20'h0a970: out <= 12'hf76;
      20'h0a971: out <= 12'hf76;
      20'h0a972: out <= 12'hf76;
      20'h0a973: out <= 12'hf76;
      20'h0a974: out <= 12'hf76;
      20'h0a975: out <= 12'hf76;
      20'h0a976: out <= 12'hf76;
      20'h0a977: out <= 12'hf76;
      20'h0a978: out <= 12'hfa9;
      20'h0a979: out <= 12'hfa9;
      20'h0a97a: out <= 12'hfa9;
      20'h0a97b: out <= 12'hfa9;
      20'h0a97c: out <= 12'hfa9;
      20'h0a97d: out <= 12'hfa9;
      20'h0a97e: out <= 12'hfa9;
      20'h0a97f: out <= 12'hfa9;
      20'h0a980: out <= 12'h000;
      20'h0a981: out <= 12'h000;
      20'h0a982: out <= 12'h000;
      20'h0a983: out <= 12'h000;
      20'h0a984: out <= 12'h000;
      20'h0a985: out <= 12'h000;
      20'h0a986: out <= 12'h000;
      20'h0a987: out <= 12'h000;
      20'h0a988: out <= 12'h088;
      20'h0a989: out <= 12'h088;
      20'h0a98a: out <= 12'h088;
      20'h0a98b: out <= 12'h088;
      20'h0a98c: out <= 12'h088;
      20'h0a98d: out <= 12'h088;
      20'h0a98e: out <= 12'h088;
      20'h0a98f: out <= 12'h088;
      20'h0a990: out <= 12'h088;
      20'h0a991: out <= 12'h088;
      20'h0a992: out <= 12'h088;
      20'h0a993: out <= 12'h088;
      20'h0a994: out <= 12'h088;
      20'h0a995: out <= 12'h088;
      20'h0a996: out <= 12'h088;
      20'h0a997: out <= 12'h088;
      20'h0a998: out <= 12'h088;
      20'h0a999: out <= 12'h088;
      20'h0a99a: out <= 12'h088;
      20'h0a99b: out <= 12'h088;
      20'h0a99c: out <= 12'h088;
      20'h0a99d: out <= 12'h088;
      20'h0a99e: out <= 12'h088;
      20'h0a99f: out <= 12'h088;
      20'h0a9a0: out <= 12'h088;
      20'h0a9a1: out <= 12'h088;
      20'h0a9a2: out <= 12'h088;
      20'h0a9a3: out <= 12'h088;
      20'h0a9a4: out <= 12'h088;
      20'h0a9a5: out <= 12'h088;
      20'h0a9a6: out <= 12'h088;
      20'h0a9a7: out <= 12'h088;
      20'h0a9a8: out <= 12'h088;
      20'h0a9a9: out <= 12'h088;
      20'h0a9aa: out <= 12'h088;
      20'h0a9ab: out <= 12'h088;
      20'h0a9ac: out <= 12'h088;
      20'h0a9ad: out <= 12'h088;
      20'h0a9ae: out <= 12'h088;
      20'h0a9af: out <= 12'h088;
      20'h0a9b0: out <= 12'h088;
      20'h0a9b1: out <= 12'h088;
      20'h0a9b2: out <= 12'h088;
      20'h0a9b3: out <= 12'h088;
      20'h0a9b4: out <= 12'h088;
      20'h0a9b5: out <= 12'h088;
      20'h0a9b6: out <= 12'h088;
      20'h0a9b7: out <= 12'h088;
      20'h0a9b8: out <= 12'h088;
      20'h0a9b9: out <= 12'h088;
      20'h0a9ba: out <= 12'h088;
      20'h0a9bb: out <= 12'h088;
      20'h0a9bc: out <= 12'h088;
      20'h0a9bd: out <= 12'h088;
      20'h0a9be: out <= 12'h088;
      20'h0a9bf: out <= 12'h088;
      20'h0a9c0: out <= 12'h088;
      20'h0a9c1: out <= 12'h088;
      20'h0a9c2: out <= 12'h088;
      20'h0a9c3: out <= 12'h088;
      20'h0a9c4: out <= 12'h088;
      20'h0a9c5: out <= 12'h088;
      20'h0a9c6: out <= 12'h088;
      20'h0a9c7: out <= 12'h088;
      20'h0a9c8: out <= 12'h088;
      20'h0a9c9: out <= 12'h088;
      20'h0a9ca: out <= 12'h088;
      20'h0a9cb: out <= 12'h088;
      20'h0a9cc: out <= 12'h088;
      20'h0a9cd: out <= 12'h088;
      20'h0a9ce: out <= 12'h088;
      20'h0a9cf: out <= 12'h088;
      20'h0a9d0: out <= 12'h088;
      20'h0a9d1: out <= 12'h088;
      20'h0a9d2: out <= 12'h088;
      20'h0a9d3: out <= 12'h088;
      20'h0a9d4: out <= 12'h088;
      20'h0a9d5: out <= 12'h088;
      20'h0a9d6: out <= 12'h088;
      20'h0a9d7: out <= 12'h088;
      20'h0a9d8: out <= 12'h088;
      20'h0a9d9: out <= 12'h088;
      20'h0a9da: out <= 12'h088;
      20'h0a9db: out <= 12'h088;
      20'h0a9dc: out <= 12'h088;
      20'h0a9dd: out <= 12'h088;
      20'h0a9de: out <= 12'h088;
      20'h0a9df: out <= 12'h088;
      20'h0a9e0: out <= 12'h088;
      20'h0a9e1: out <= 12'h088;
      20'h0a9e2: out <= 12'h088;
      20'h0a9e3: out <= 12'h088;
      20'h0a9e4: out <= 12'h088;
      20'h0a9e5: out <= 12'h088;
      20'h0a9e6: out <= 12'h088;
      20'h0a9e7: out <= 12'h088;
      20'h0a9e8: out <= 12'h088;
      20'h0a9e9: out <= 12'h088;
      20'h0a9ea: out <= 12'h088;
      20'h0a9eb: out <= 12'h088;
      20'h0a9ec: out <= 12'h088;
      20'h0a9ed: out <= 12'h088;
      20'h0a9ee: out <= 12'h088;
      20'h0a9ef: out <= 12'h088;
      20'h0a9f0: out <= 12'h088;
      20'h0a9f1: out <= 12'hbb0;
      20'h0a9f2: out <= 12'h660;
      20'h0a9f3: out <= 12'h660;
      20'h0a9f4: out <= 12'h660;
      20'h0a9f5: out <= 12'h660;
      20'h0a9f6: out <= 12'h660;
      20'h0a9f7: out <= 12'h660;
      20'h0a9f8: out <= 12'h222;
      20'h0a9f9: out <= 12'h660;
      20'h0a9fa: out <= 12'h660;
      20'h0a9fb: out <= 12'h660;
      20'h0a9fc: out <= 12'hbb0;
      20'h0a9fd: out <= 12'hee9;
      20'h0a9fe: out <= 12'hee9;
      20'h0a9ff: out <= 12'h660;
      20'h0aa00: out <= 12'hee9;
      20'h0aa01: out <= 12'hbb0;
      20'h0aa02: out <= 12'h660;
      20'h0aa03: out <= 12'h660;
      20'h0aa04: out <= 12'h660;
      20'h0aa05: out <= 12'h660;
      20'h0aa06: out <= 12'hee9;
      20'h0aa07: out <= 12'h660;
      20'h0aa08: out <= 12'h603;
      20'h0aa09: out <= 12'h603;
      20'h0aa0a: out <= 12'h603;
      20'h0aa0b: out <= 12'h603;
      20'h0aa0c: out <= 12'hbbb;
      20'h0aa0d: out <= 12'hbbb;
      20'h0aa0e: out <= 12'h000;
      20'h0aa0f: out <= 12'hbbb;
      20'h0aa10: out <= 12'h000;
      20'h0aa11: out <= 12'hbbb;
      20'h0aa12: out <= 12'hbbb;
      20'h0aa13: out <= 12'h000;
      20'h0aa14: out <= 12'h000;
      20'h0aa15: out <= 12'h000;
      20'h0aa16: out <= 12'h000;
      20'h0aa17: out <= 12'hbbb;
      20'h0aa18: out <= 12'hbbb;
      20'h0aa19: out <= 12'h000;
      20'h0aa1a: out <= 12'h000;
      20'h0aa1b: out <= 12'h000;
      20'h0aa1c: out <= 12'h000;
      20'h0aa1d: out <= 12'h000;
      20'h0aa1e: out <= 12'h000;
      20'h0aa1f: out <= 12'hbbb;
      20'h0aa20: out <= 12'hbbb;
      20'h0aa21: out <= 12'hbbb;
      20'h0aa22: out <= 12'h000;
      20'h0aa23: out <= 12'h000;
      20'h0aa24: out <= 12'h000;
      20'h0aa25: out <= 12'h000;
      20'h0aa26: out <= 12'hbbb;
      20'h0aa27: out <= 12'hbbb;
      20'h0aa28: out <= 12'hbbb;
      20'h0aa29: out <= 12'hbbb;
      20'h0aa2a: out <= 12'h000;
      20'h0aa2b: out <= 12'h000;
      20'h0aa2c: out <= 12'hbbb;
      20'h0aa2d: out <= 12'hbbb;
      20'h0aa2e: out <= 12'h000;
      20'h0aa2f: out <= 12'h000;
      20'h0aa30: out <= 12'hbbb;
      20'h0aa31: out <= 12'hbbb;
      20'h0aa32: out <= 12'h000;
      20'h0aa33: out <= 12'h000;
      20'h0aa34: out <= 12'h000;
      20'h0aa35: out <= 12'h000;
      20'h0aa36: out <= 12'h000;
      20'h0aa37: out <= 12'h000;
      20'h0aa38: out <= 12'h000;
      20'h0aa39: out <= 12'hbbb;
      20'h0aa3a: out <= 12'hbbb;
      20'h0aa3b: out <= 12'h000;
      20'h0aa3c: out <= 12'hbbb;
      20'h0aa3d: out <= 12'hbbb;
      20'h0aa3e: out <= 12'hbbb;
      20'h0aa3f: out <= 12'hbbb;
      20'h0aa40: out <= 12'hbbb;
      20'h0aa41: out <= 12'hbbb;
      20'h0aa42: out <= 12'h000;
      20'h0aa43: out <= 12'h000;
      20'h0aa44: out <= 12'h000;
      20'h0aa45: out <= 12'h000;
      20'h0aa46: out <= 12'h000;
      20'h0aa47: out <= 12'hbbb;
      20'h0aa48: out <= 12'hbbb;
      20'h0aa49: out <= 12'h000;
      20'h0aa4a: out <= 12'h000;
      20'h0aa4b: out <= 12'h000;
      20'h0aa4c: out <= 12'h000;
      20'h0aa4d: out <= 12'hbbb;
      20'h0aa4e: out <= 12'hbbb;
      20'h0aa4f: out <= 12'hbbb;
      20'h0aa50: out <= 12'hbbb;
      20'h0aa51: out <= 12'hbbb;
      20'h0aa52: out <= 12'h000;
      20'h0aa53: out <= 12'h000;
      20'h0aa54: out <= 12'h000;
      20'h0aa55: out <= 12'hbbb;
      20'h0aa56: out <= 12'hbbb;
      20'h0aa57: out <= 12'hbbb;
      20'h0aa58: out <= 12'hbbb;
      20'h0aa59: out <= 12'hbbb;
      20'h0aa5a: out <= 12'hbbb;
      20'h0aa5b: out <= 12'h000;
      20'h0aa5c: out <= 12'h603;
      20'h0aa5d: out <= 12'h603;
      20'h0aa5e: out <= 12'h603;
      20'h0aa5f: out <= 12'h603;
      20'h0aa60: out <= 12'hee9;
      20'h0aa61: out <= 12'hf87;
      20'h0aa62: out <= 12'hee9;
      20'h0aa63: out <= 12'hf87;
      20'h0aa64: out <= 12'hf87;
      20'h0aa65: out <= 12'hb27;
      20'h0aa66: out <= 12'hf87;
      20'h0aa67: out <= 12'hb27;
      20'h0aa68: out <= 12'h000;
      20'h0aa69: out <= 12'h000;
      20'h0aa6a: out <= 12'h000;
      20'h0aa6b: out <= 12'h000;
      20'h0aa6c: out <= 12'h000;
      20'h0aa6d: out <= 12'h000;
      20'h0aa6e: out <= 12'h000;
      20'h0aa6f: out <= 12'h000;
      20'h0aa70: out <= 12'hfa9;
      20'h0aa71: out <= 12'hfa9;
      20'h0aa72: out <= 12'hfa9;
      20'h0aa73: out <= 12'hfa9;
      20'h0aa74: out <= 12'hfa9;
      20'h0aa75: out <= 12'hfa9;
      20'h0aa76: out <= 12'hfa9;
      20'h0aa77: out <= 12'hfa9;
      20'h0aa78: out <= 12'hf76;
      20'h0aa79: out <= 12'hf76;
      20'h0aa7a: out <= 12'hf76;
      20'h0aa7b: out <= 12'hf76;
      20'h0aa7c: out <= 12'hf76;
      20'h0aa7d: out <= 12'hf76;
      20'h0aa7e: out <= 12'hf76;
      20'h0aa7f: out <= 12'hf76;
      20'h0aa80: out <= 12'hfa9;
      20'h0aa81: out <= 12'hfa9;
      20'h0aa82: out <= 12'hfa9;
      20'h0aa83: out <= 12'hfa9;
      20'h0aa84: out <= 12'hfa9;
      20'h0aa85: out <= 12'hfa9;
      20'h0aa86: out <= 12'hfa9;
      20'h0aa87: out <= 12'hfa9;
      20'h0aa88: out <= 12'hf76;
      20'h0aa89: out <= 12'hf76;
      20'h0aa8a: out <= 12'hf76;
      20'h0aa8b: out <= 12'hf76;
      20'h0aa8c: out <= 12'hf76;
      20'h0aa8d: out <= 12'hf76;
      20'h0aa8e: out <= 12'hf76;
      20'h0aa8f: out <= 12'hf76;
      20'h0aa90: out <= 12'hfa9;
      20'h0aa91: out <= 12'hfa9;
      20'h0aa92: out <= 12'hfa9;
      20'h0aa93: out <= 12'hfa9;
      20'h0aa94: out <= 12'hfa9;
      20'h0aa95: out <= 12'hfa9;
      20'h0aa96: out <= 12'hfa9;
      20'h0aa97: out <= 12'hfa9;
      20'h0aa98: out <= 12'h000;
      20'h0aa99: out <= 12'h000;
      20'h0aa9a: out <= 12'h000;
      20'h0aa9b: out <= 12'h000;
      20'h0aa9c: out <= 12'h000;
      20'h0aa9d: out <= 12'h000;
      20'h0aa9e: out <= 12'h000;
      20'h0aa9f: out <= 12'h000;
      20'h0aaa0: out <= 12'h088;
      20'h0aaa1: out <= 12'h088;
      20'h0aaa2: out <= 12'h088;
      20'h0aaa3: out <= 12'h088;
      20'h0aaa4: out <= 12'h088;
      20'h0aaa5: out <= 12'h088;
      20'h0aaa6: out <= 12'h088;
      20'h0aaa7: out <= 12'h088;
      20'h0aaa8: out <= 12'h088;
      20'h0aaa9: out <= 12'h088;
      20'h0aaaa: out <= 12'h088;
      20'h0aaab: out <= 12'h088;
      20'h0aaac: out <= 12'h088;
      20'h0aaad: out <= 12'h088;
      20'h0aaae: out <= 12'h088;
      20'h0aaaf: out <= 12'h088;
      20'h0aab0: out <= 12'h088;
      20'h0aab1: out <= 12'h088;
      20'h0aab2: out <= 12'h088;
      20'h0aab3: out <= 12'h088;
      20'h0aab4: out <= 12'h088;
      20'h0aab5: out <= 12'h088;
      20'h0aab6: out <= 12'h088;
      20'h0aab7: out <= 12'h088;
      20'h0aab8: out <= 12'h088;
      20'h0aab9: out <= 12'h088;
      20'h0aaba: out <= 12'h088;
      20'h0aabb: out <= 12'h088;
      20'h0aabc: out <= 12'h088;
      20'h0aabd: out <= 12'h088;
      20'h0aabe: out <= 12'h088;
      20'h0aabf: out <= 12'h088;
      20'h0aac0: out <= 12'h088;
      20'h0aac1: out <= 12'h088;
      20'h0aac2: out <= 12'h088;
      20'h0aac3: out <= 12'h088;
      20'h0aac4: out <= 12'h088;
      20'h0aac5: out <= 12'h088;
      20'h0aac6: out <= 12'h088;
      20'h0aac7: out <= 12'h088;
      20'h0aac8: out <= 12'h088;
      20'h0aac9: out <= 12'h088;
      20'h0aaca: out <= 12'h088;
      20'h0aacb: out <= 12'h088;
      20'h0aacc: out <= 12'h088;
      20'h0aacd: out <= 12'h088;
      20'h0aace: out <= 12'h088;
      20'h0aacf: out <= 12'h088;
      20'h0aad0: out <= 12'h088;
      20'h0aad1: out <= 12'h088;
      20'h0aad2: out <= 12'h088;
      20'h0aad3: out <= 12'h088;
      20'h0aad4: out <= 12'h088;
      20'h0aad5: out <= 12'h088;
      20'h0aad6: out <= 12'h088;
      20'h0aad7: out <= 12'h088;
      20'h0aad8: out <= 12'h088;
      20'h0aad9: out <= 12'h088;
      20'h0aada: out <= 12'h088;
      20'h0aadb: out <= 12'h088;
      20'h0aadc: out <= 12'h088;
      20'h0aadd: out <= 12'h088;
      20'h0aade: out <= 12'h088;
      20'h0aadf: out <= 12'h088;
      20'h0aae0: out <= 12'h088;
      20'h0aae1: out <= 12'h088;
      20'h0aae2: out <= 12'h088;
      20'h0aae3: out <= 12'h088;
      20'h0aae4: out <= 12'h088;
      20'h0aae5: out <= 12'h088;
      20'h0aae6: out <= 12'h088;
      20'h0aae7: out <= 12'h088;
      20'h0aae8: out <= 12'h088;
      20'h0aae9: out <= 12'h088;
      20'h0aaea: out <= 12'h088;
      20'h0aaeb: out <= 12'h088;
      20'h0aaec: out <= 12'h088;
      20'h0aaed: out <= 12'h088;
      20'h0aaee: out <= 12'h088;
      20'h0aaef: out <= 12'h088;
      20'h0aaf0: out <= 12'h088;
      20'h0aaf1: out <= 12'h088;
      20'h0aaf2: out <= 12'h088;
      20'h0aaf3: out <= 12'h088;
      20'h0aaf4: out <= 12'h088;
      20'h0aaf5: out <= 12'h088;
      20'h0aaf6: out <= 12'h088;
      20'h0aaf7: out <= 12'h088;
      20'h0aaf8: out <= 12'h088;
      20'h0aaf9: out <= 12'h088;
      20'h0aafa: out <= 12'h088;
      20'h0aafb: out <= 12'h088;
      20'h0aafc: out <= 12'h088;
      20'h0aafd: out <= 12'h088;
      20'h0aafe: out <= 12'h088;
      20'h0aaff: out <= 12'h088;
      20'h0ab00: out <= 12'h088;
      20'h0ab01: out <= 12'h088;
      20'h0ab02: out <= 12'h088;
      20'h0ab03: out <= 12'h088;
      20'h0ab04: out <= 12'h088;
      20'h0ab05: out <= 12'h088;
      20'h0ab06: out <= 12'h088;
      20'h0ab07: out <= 12'h088;
      20'h0ab08: out <= 12'h088;
      20'h0ab09: out <= 12'hbb0;
      20'h0ab0a: out <= 12'h660;
      20'h0ab0b: out <= 12'h660;
      20'h0ab0c: out <= 12'h660;
      20'h0ab0d: out <= 12'hbb0;
      20'h0ab0e: out <= 12'hee9;
      20'h0ab0f: out <= 12'h660;
      20'h0ab10: out <= 12'h222;
      20'h0ab11: out <= 12'h660;
      20'h0ab12: out <= 12'hee9;
      20'h0ab13: out <= 12'hbb0;
      20'h0ab14: out <= 12'hbb0;
      20'h0ab15: out <= 12'hee9;
      20'h0ab16: out <= 12'hee9;
      20'h0ab17: out <= 12'h660;
      20'h0ab18: out <= 12'hee9;
      20'h0ab19: out <= 12'hbb0;
      20'h0ab1a: out <= 12'h660;
      20'h0ab1b: out <= 12'h660;
      20'h0ab1c: out <= 12'h660;
      20'h0ab1d: out <= 12'hbb0;
      20'h0ab1e: out <= 12'h660;
      20'h0ab1f: out <= 12'h660;
      20'h0ab20: out <= 12'h603;
      20'h0ab21: out <= 12'h603;
      20'h0ab22: out <= 12'h603;
      20'h0ab23: out <= 12'h603;
      20'h0ab24: out <= 12'hbbb;
      20'h0ab25: out <= 12'hbbb;
      20'h0ab26: out <= 12'hbbb;
      20'h0ab27: out <= 12'h000;
      20'h0ab28: out <= 12'h000;
      20'h0ab29: out <= 12'hbbb;
      20'h0ab2a: out <= 12'hbbb;
      20'h0ab2b: out <= 12'h000;
      20'h0ab2c: out <= 12'h000;
      20'h0ab2d: out <= 12'h000;
      20'h0ab2e: out <= 12'h000;
      20'h0ab2f: out <= 12'hbbb;
      20'h0ab30: out <= 12'hbbb;
      20'h0ab31: out <= 12'h000;
      20'h0ab32: out <= 12'h000;
      20'h0ab33: out <= 12'h000;
      20'h0ab34: out <= 12'h000;
      20'h0ab35: out <= 12'hbbb;
      20'h0ab36: out <= 12'hbbb;
      20'h0ab37: out <= 12'hbbb;
      20'h0ab38: out <= 12'h000;
      20'h0ab39: out <= 12'h000;
      20'h0ab3a: out <= 12'h000;
      20'h0ab3b: out <= 12'h000;
      20'h0ab3c: out <= 12'h000;
      20'h0ab3d: out <= 12'h000;
      20'h0ab3e: out <= 12'h000;
      20'h0ab3f: out <= 12'h000;
      20'h0ab40: out <= 12'h000;
      20'h0ab41: out <= 12'hbbb;
      20'h0ab42: out <= 12'hbbb;
      20'h0ab43: out <= 12'h000;
      20'h0ab44: out <= 12'hbbb;
      20'h0ab45: out <= 12'hbbb;
      20'h0ab46: out <= 12'hbbb;
      20'h0ab47: out <= 12'hbbb;
      20'h0ab48: out <= 12'hbbb;
      20'h0ab49: out <= 12'hbbb;
      20'h0ab4a: out <= 12'hbbb;
      20'h0ab4b: out <= 12'h000;
      20'h0ab4c: out <= 12'h000;
      20'h0ab4d: out <= 12'h000;
      20'h0ab4e: out <= 12'h000;
      20'h0ab4f: out <= 12'h000;
      20'h0ab50: out <= 12'h000;
      20'h0ab51: out <= 12'hbbb;
      20'h0ab52: out <= 12'hbbb;
      20'h0ab53: out <= 12'h000;
      20'h0ab54: out <= 12'hbbb;
      20'h0ab55: out <= 12'hbbb;
      20'h0ab56: out <= 12'h000;
      20'h0ab57: out <= 12'h000;
      20'h0ab58: out <= 12'h000;
      20'h0ab59: out <= 12'hbbb;
      20'h0ab5a: out <= 12'hbbb;
      20'h0ab5b: out <= 12'h000;
      20'h0ab5c: out <= 12'h000;
      20'h0ab5d: out <= 12'h000;
      20'h0ab5e: out <= 12'hbbb;
      20'h0ab5f: out <= 12'hbbb;
      20'h0ab60: out <= 12'h000;
      20'h0ab61: out <= 12'h000;
      20'h0ab62: out <= 12'h000;
      20'h0ab63: out <= 12'h000;
      20'h0ab64: out <= 12'hbbb;
      20'h0ab65: out <= 12'hbbb;
      20'h0ab66: out <= 12'h000;
      20'h0ab67: out <= 12'h000;
      20'h0ab68: out <= 12'h000;
      20'h0ab69: out <= 12'hbbb;
      20'h0ab6a: out <= 12'hbbb;
      20'h0ab6b: out <= 12'h000;
      20'h0ab6c: out <= 12'h000;
      20'h0ab6d: out <= 12'h000;
      20'h0ab6e: out <= 12'h000;
      20'h0ab6f: out <= 12'h000;
      20'h0ab70: out <= 12'h000;
      20'h0ab71: out <= 12'hbbb;
      20'h0ab72: out <= 12'hbbb;
      20'h0ab73: out <= 12'h000;
      20'h0ab74: out <= 12'h603;
      20'h0ab75: out <= 12'h603;
      20'h0ab76: out <= 12'h603;
      20'h0ab77: out <= 12'h603;
      20'h0ab78: out <= 12'hee9;
      20'h0ab79: out <= 12'hf87;
      20'h0ab7a: out <= 12'hee9;
      20'h0ab7b: out <= 12'hf87;
      20'h0ab7c: out <= 12'hf87;
      20'h0ab7d: out <= 12'hb27;
      20'h0ab7e: out <= 12'hf87;
      20'h0ab7f: out <= 12'hb27;
      20'h0ab80: out <= 12'h000;
      20'h0ab81: out <= 12'h000;
      20'h0ab82: out <= 12'h000;
      20'h0ab83: out <= 12'h000;
      20'h0ab84: out <= 12'h000;
      20'h0ab85: out <= 12'h000;
      20'h0ab86: out <= 12'h000;
      20'h0ab87: out <= 12'h000;
      20'h0ab88: out <= 12'hfa9;
      20'h0ab89: out <= 12'hfa9;
      20'h0ab8a: out <= 12'hfa9;
      20'h0ab8b: out <= 12'hfa9;
      20'h0ab8c: out <= 12'hfa9;
      20'h0ab8d: out <= 12'hfa9;
      20'h0ab8e: out <= 12'hfa9;
      20'h0ab8f: out <= 12'hfa9;
      20'h0ab90: out <= 12'hf76;
      20'h0ab91: out <= 12'hf76;
      20'h0ab92: out <= 12'hf76;
      20'h0ab93: out <= 12'hf76;
      20'h0ab94: out <= 12'hf76;
      20'h0ab95: out <= 12'hf76;
      20'h0ab96: out <= 12'hf76;
      20'h0ab97: out <= 12'hf76;
      20'h0ab98: out <= 12'hfa9;
      20'h0ab99: out <= 12'hfa9;
      20'h0ab9a: out <= 12'hfa9;
      20'h0ab9b: out <= 12'hfa9;
      20'h0ab9c: out <= 12'hfa9;
      20'h0ab9d: out <= 12'hfa9;
      20'h0ab9e: out <= 12'hfa9;
      20'h0ab9f: out <= 12'hfa9;
      20'h0aba0: out <= 12'hf76;
      20'h0aba1: out <= 12'hf76;
      20'h0aba2: out <= 12'hf76;
      20'h0aba3: out <= 12'hf76;
      20'h0aba4: out <= 12'hf76;
      20'h0aba5: out <= 12'hf76;
      20'h0aba6: out <= 12'hf76;
      20'h0aba7: out <= 12'hf76;
      20'h0aba8: out <= 12'hfa9;
      20'h0aba9: out <= 12'hfa9;
      20'h0abaa: out <= 12'hfa9;
      20'h0abab: out <= 12'hfa9;
      20'h0abac: out <= 12'hfa9;
      20'h0abad: out <= 12'hfa9;
      20'h0abae: out <= 12'hfa9;
      20'h0abaf: out <= 12'hfa9;
      20'h0abb0: out <= 12'h000;
      20'h0abb1: out <= 12'h000;
      20'h0abb2: out <= 12'h000;
      20'h0abb3: out <= 12'h000;
      20'h0abb4: out <= 12'h000;
      20'h0abb5: out <= 12'h000;
      20'h0abb6: out <= 12'h000;
      20'h0abb7: out <= 12'h000;
      20'h0abb8: out <= 12'h088;
      20'h0abb9: out <= 12'h088;
      20'h0abba: out <= 12'h088;
      20'h0abbb: out <= 12'h088;
      20'h0abbc: out <= 12'h088;
      20'h0abbd: out <= 12'h088;
      20'h0abbe: out <= 12'h088;
      20'h0abbf: out <= 12'h088;
      20'h0abc0: out <= 12'h088;
      20'h0abc1: out <= 12'h088;
      20'h0abc2: out <= 12'h088;
      20'h0abc3: out <= 12'h088;
      20'h0abc4: out <= 12'h088;
      20'h0abc5: out <= 12'h088;
      20'h0abc6: out <= 12'h088;
      20'h0abc7: out <= 12'h088;
      20'h0abc8: out <= 12'h088;
      20'h0abc9: out <= 12'h088;
      20'h0abca: out <= 12'h088;
      20'h0abcb: out <= 12'h088;
      20'h0abcc: out <= 12'h088;
      20'h0abcd: out <= 12'h088;
      20'h0abce: out <= 12'h088;
      20'h0abcf: out <= 12'h088;
      20'h0abd0: out <= 12'h088;
      20'h0abd1: out <= 12'h088;
      20'h0abd2: out <= 12'h088;
      20'h0abd3: out <= 12'h088;
      20'h0abd4: out <= 12'h088;
      20'h0abd5: out <= 12'h088;
      20'h0abd6: out <= 12'h088;
      20'h0abd7: out <= 12'h088;
      20'h0abd8: out <= 12'h088;
      20'h0abd9: out <= 12'h088;
      20'h0abda: out <= 12'h088;
      20'h0abdb: out <= 12'h088;
      20'h0abdc: out <= 12'h088;
      20'h0abdd: out <= 12'h088;
      20'h0abde: out <= 12'h088;
      20'h0abdf: out <= 12'h088;
      20'h0abe0: out <= 12'h088;
      20'h0abe1: out <= 12'h088;
      20'h0abe2: out <= 12'h088;
      20'h0abe3: out <= 12'h088;
      20'h0abe4: out <= 12'h088;
      20'h0abe5: out <= 12'h088;
      20'h0abe6: out <= 12'h088;
      20'h0abe7: out <= 12'h088;
      20'h0abe8: out <= 12'h088;
      20'h0abe9: out <= 12'h088;
      20'h0abea: out <= 12'h088;
      20'h0abeb: out <= 12'h088;
      20'h0abec: out <= 12'h088;
      20'h0abed: out <= 12'h088;
      20'h0abee: out <= 12'h088;
      20'h0abef: out <= 12'h088;
      20'h0abf0: out <= 12'h088;
      20'h0abf1: out <= 12'h088;
      20'h0abf2: out <= 12'h088;
      20'h0abf3: out <= 12'h088;
      20'h0abf4: out <= 12'h088;
      20'h0abf5: out <= 12'h088;
      20'h0abf6: out <= 12'h088;
      20'h0abf7: out <= 12'h088;
      20'h0abf8: out <= 12'h088;
      20'h0abf9: out <= 12'h088;
      20'h0abfa: out <= 12'h088;
      20'h0abfb: out <= 12'h088;
      20'h0abfc: out <= 12'h088;
      20'h0abfd: out <= 12'h088;
      20'h0abfe: out <= 12'h088;
      20'h0abff: out <= 12'h088;
      20'h0ac00: out <= 12'h088;
      20'h0ac01: out <= 12'h088;
      20'h0ac02: out <= 12'h088;
      20'h0ac03: out <= 12'h088;
      20'h0ac04: out <= 12'h088;
      20'h0ac05: out <= 12'h088;
      20'h0ac06: out <= 12'h088;
      20'h0ac07: out <= 12'h088;
      20'h0ac08: out <= 12'h088;
      20'h0ac09: out <= 12'h088;
      20'h0ac0a: out <= 12'h088;
      20'h0ac0b: out <= 12'h088;
      20'h0ac0c: out <= 12'h088;
      20'h0ac0d: out <= 12'h088;
      20'h0ac0e: out <= 12'h088;
      20'h0ac0f: out <= 12'h088;
      20'h0ac10: out <= 12'h088;
      20'h0ac11: out <= 12'h088;
      20'h0ac12: out <= 12'h088;
      20'h0ac13: out <= 12'h088;
      20'h0ac14: out <= 12'h088;
      20'h0ac15: out <= 12'h088;
      20'h0ac16: out <= 12'h088;
      20'h0ac17: out <= 12'h088;
      20'h0ac18: out <= 12'h088;
      20'h0ac19: out <= 12'h088;
      20'h0ac1a: out <= 12'h088;
      20'h0ac1b: out <= 12'h088;
      20'h0ac1c: out <= 12'h088;
      20'h0ac1d: out <= 12'h088;
      20'h0ac1e: out <= 12'h088;
      20'h0ac1f: out <= 12'h088;
      20'h0ac20: out <= 12'h088;
      20'h0ac21: out <= 12'hbb0;
      20'h0ac22: out <= 12'h660;
      20'h0ac23: out <= 12'h660;
      20'h0ac24: out <= 12'h660;
      20'h0ac25: out <= 12'hbb0;
      20'h0ac26: out <= 12'h660;
      20'h0ac27: out <= 12'h660;
      20'h0ac28: out <= 12'h222;
      20'h0ac29: out <= 12'h660;
      20'h0ac2a: out <= 12'h660;
      20'h0ac2b: out <= 12'hbb0;
      20'h0ac2c: out <= 12'hbb0;
      20'h0ac2d: out <= 12'hee9;
      20'h0ac2e: out <= 12'hee9;
      20'h0ac2f: out <= 12'h660;
      20'h0ac30: out <= 12'hee9;
      20'h0ac31: out <= 12'hbb0;
      20'h0ac32: out <= 12'h660;
      20'h0ac33: out <= 12'h660;
      20'h0ac34: out <= 12'h660;
      20'h0ac35: out <= 12'hbb0;
      20'h0ac36: out <= 12'hee9;
      20'h0ac37: out <= 12'h660;
      20'h0ac38: out <= 12'h603;
      20'h0ac39: out <= 12'h603;
      20'h0ac3a: out <= 12'h603;
      20'h0ac3b: out <= 12'h603;
      20'h0ac3c: out <= 12'hbbb;
      20'h0ac3d: out <= 12'hbbb;
      20'h0ac3e: out <= 12'h000;
      20'h0ac3f: out <= 12'h000;
      20'h0ac40: out <= 12'h000;
      20'h0ac41: out <= 12'hbbb;
      20'h0ac42: out <= 12'hbbb;
      20'h0ac43: out <= 12'h000;
      20'h0ac44: out <= 12'h000;
      20'h0ac45: out <= 12'h000;
      20'h0ac46: out <= 12'h000;
      20'h0ac47: out <= 12'hbbb;
      20'h0ac48: out <= 12'hbbb;
      20'h0ac49: out <= 12'h000;
      20'h0ac4a: out <= 12'h000;
      20'h0ac4b: out <= 12'h000;
      20'h0ac4c: out <= 12'hbbb;
      20'h0ac4d: out <= 12'hbbb;
      20'h0ac4e: out <= 12'h000;
      20'h0ac4f: out <= 12'h000;
      20'h0ac50: out <= 12'h000;
      20'h0ac51: out <= 12'h000;
      20'h0ac52: out <= 12'h000;
      20'h0ac53: out <= 12'h000;
      20'h0ac54: out <= 12'hbbb;
      20'h0ac55: out <= 12'hbbb;
      20'h0ac56: out <= 12'h000;
      20'h0ac57: out <= 12'h000;
      20'h0ac58: out <= 12'h000;
      20'h0ac59: out <= 12'hbbb;
      20'h0ac5a: out <= 12'hbbb;
      20'h0ac5b: out <= 12'h000;
      20'h0ac5c: out <= 12'h000;
      20'h0ac5d: out <= 12'h000;
      20'h0ac5e: out <= 12'h000;
      20'h0ac5f: out <= 12'h000;
      20'h0ac60: out <= 12'hbbb;
      20'h0ac61: out <= 12'hbbb;
      20'h0ac62: out <= 12'h000;
      20'h0ac63: out <= 12'h000;
      20'h0ac64: out <= 12'hbbb;
      20'h0ac65: out <= 12'hbbb;
      20'h0ac66: out <= 12'h000;
      20'h0ac67: out <= 12'h000;
      20'h0ac68: out <= 12'h000;
      20'h0ac69: out <= 12'hbbb;
      20'h0ac6a: out <= 12'hbbb;
      20'h0ac6b: out <= 12'h000;
      20'h0ac6c: out <= 12'hbbb;
      20'h0ac6d: out <= 12'hbbb;
      20'h0ac6e: out <= 12'h000;
      20'h0ac6f: out <= 12'h000;
      20'h0ac70: out <= 12'h000;
      20'h0ac71: out <= 12'hbbb;
      20'h0ac72: out <= 12'hbbb;
      20'h0ac73: out <= 12'h000;
      20'h0ac74: out <= 12'h000;
      20'h0ac75: out <= 12'h000;
      20'h0ac76: out <= 12'hbbb;
      20'h0ac77: out <= 12'hbbb;
      20'h0ac78: out <= 12'h000;
      20'h0ac79: out <= 12'h000;
      20'h0ac7a: out <= 12'h000;
      20'h0ac7b: out <= 12'h000;
      20'h0ac7c: out <= 12'hbbb;
      20'h0ac7d: out <= 12'hbbb;
      20'h0ac7e: out <= 12'h000;
      20'h0ac7f: out <= 12'h000;
      20'h0ac80: out <= 12'h000;
      20'h0ac81: out <= 12'hbbb;
      20'h0ac82: out <= 12'hbbb;
      20'h0ac83: out <= 12'h000;
      20'h0ac84: out <= 12'h000;
      20'h0ac85: out <= 12'h000;
      20'h0ac86: out <= 12'h000;
      20'h0ac87: out <= 12'h000;
      20'h0ac88: out <= 12'hbbb;
      20'h0ac89: out <= 12'hbbb;
      20'h0ac8a: out <= 12'h000;
      20'h0ac8b: out <= 12'h000;
      20'h0ac8c: out <= 12'h603;
      20'h0ac8d: out <= 12'h603;
      20'h0ac8e: out <= 12'h603;
      20'h0ac8f: out <= 12'h603;
      20'h0ac90: out <= 12'hee9;
      20'h0ac91: out <= 12'hf87;
      20'h0ac92: out <= 12'hee9;
      20'h0ac93: out <= 12'hb27;
      20'h0ac94: out <= 12'hb27;
      20'h0ac95: out <= 12'hb27;
      20'h0ac96: out <= 12'hf87;
      20'h0ac97: out <= 12'hb27;
      20'h0ac98: out <= 12'h000;
      20'h0ac99: out <= 12'h000;
      20'h0ac9a: out <= 12'h000;
      20'h0ac9b: out <= 12'h000;
      20'h0ac9c: out <= 12'h000;
      20'h0ac9d: out <= 12'h000;
      20'h0ac9e: out <= 12'h000;
      20'h0ac9f: out <= 12'h000;
      20'h0aca0: out <= 12'hfa9;
      20'h0aca1: out <= 12'hfa9;
      20'h0aca2: out <= 12'hfa9;
      20'h0aca3: out <= 12'hfa9;
      20'h0aca4: out <= 12'hfa9;
      20'h0aca5: out <= 12'hfa9;
      20'h0aca6: out <= 12'hfa9;
      20'h0aca7: out <= 12'hfa9;
      20'h0aca8: out <= 12'hf76;
      20'h0aca9: out <= 12'hf76;
      20'h0acaa: out <= 12'hf76;
      20'h0acab: out <= 12'hf76;
      20'h0acac: out <= 12'hf76;
      20'h0acad: out <= 12'hf76;
      20'h0acae: out <= 12'hf76;
      20'h0acaf: out <= 12'hf76;
      20'h0acb0: out <= 12'hfa9;
      20'h0acb1: out <= 12'hfa9;
      20'h0acb2: out <= 12'hfa9;
      20'h0acb3: out <= 12'hfa9;
      20'h0acb4: out <= 12'hfa9;
      20'h0acb5: out <= 12'hfa9;
      20'h0acb6: out <= 12'hfa9;
      20'h0acb7: out <= 12'hfa9;
      20'h0acb8: out <= 12'hf76;
      20'h0acb9: out <= 12'hf76;
      20'h0acba: out <= 12'hf76;
      20'h0acbb: out <= 12'hf76;
      20'h0acbc: out <= 12'hf76;
      20'h0acbd: out <= 12'hf76;
      20'h0acbe: out <= 12'hf76;
      20'h0acbf: out <= 12'hf76;
      20'h0acc0: out <= 12'hfa9;
      20'h0acc1: out <= 12'hfa9;
      20'h0acc2: out <= 12'hfa9;
      20'h0acc3: out <= 12'hfa9;
      20'h0acc4: out <= 12'hfa9;
      20'h0acc5: out <= 12'hfa9;
      20'h0acc6: out <= 12'hfa9;
      20'h0acc7: out <= 12'hfa9;
      20'h0acc8: out <= 12'h000;
      20'h0acc9: out <= 12'h000;
      20'h0acca: out <= 12'h000;
      20'h0accb: out <= 12'h000;
      20'h0accc: out <= 12'h000;
      20'h0accd: out <= 12'h000;
      20'h0acce: out <= 12'h000;
      20'h0accf: out <= 12'h000;
      20'h0acd0: out <= 12'h088;
      20'h0acd1: out <= 12'h088;
      20'h0acd2: out <= 12'h088;
      20'h0acd3: out <= 12'h088;
      20'h0acd4: out <= 12'h088;
      20'h0acd5: out <= 12'h088;
      20'h0acd6: out <= 12'h088;
      20'h0acd7: out <= 12'h088;
      20'h0acd8: out <= 12'h088;
      20'h0acd9: out <= 12'h088;
      20'h0acda: out <= 12'h088;
      20'h0acdb: out <= 12'h088;
      20'h0acdc: out <= 12'h088;
      20'h0acdd: out <= 12'h088;
      20'h0acde: out <= 12'h088;
      20'h0acdf: out <= 12'h088;
      20'h0ace0: out <= 12'h088;
      20'h0ace1: out <= 12'h088;
      20'h0ace2: out <= 12'h088;
      20'h0ace3: out <= 12'h088;
      20'h0ace4: out <= 12'h088;
      20'h0ace5: out <= 12'h088;
      20'h0ace6: out <= 12'h088;
      20'h0ace7: out <= 12'h088;
      20'h0ace8: out <= 12'h088;
      20'h0ace9: out <= 12'h088;
      20'h0acea: out <= 12'h088;
      20'h0aceb: out <= 12'h088;
      20'h0acec: out <= 12'h088;
      20'h0aced: out <= 12'h088;
      20'h0acee: out <= 12'h088;
      20'h0acef: out <= 12'h088;
      20'h0acf0: out <= 12'h088;
      20'h0acf1: out <= 12'h088;
      20'h0acf2: out <= 12'h088;
      20'h0acf3: out <= 12'h088;
      20'h0acf4: out <= 12'h088;
      20'h0acf5: out <= 12'h088;
      20'h0acf6: out <= 12'h088;
      20'h0acf7: out <= 12'h088;
      20'h0acf8: out <= 12'h088;
      20'h0acf9: out <= 12'h088;
      20'h0acfa: out <= 12'h088;
      20'h0acfb: out <= 12'h088;
      20'h0acfc: out <= 12'h088;
      20'h0acfd: out <= 12'h088;
      20'h0acfe: out <= 12'h088;
      20'h0acff: out <= 12'h088;
      20'h0ad00: out <= 12'h088;
      20'h0ad01: out <= 12'h088;
      20'h0ad02: out <= 12'h088;
      20'h0ad03: out <= 12'h088;
      20'h0ad04: out <= 12'h088;
      20'h0ad05: out <= 12'h088;
      20'h0ad06: out <= 12'h088;
      20'h0ad07: out <= 12'h088;
      20'h0ad08: out <= 12'h088;
      20'h0ad09: out <= 12'h088;
      20'h0ad0a: out <= 12'h088;
      20'h0ad0b: out <= 12'h088;
      20'h0ad0c: out <= 12'h088;
      20'h0ad0d: out <= 12'h088;
      20'h0ad0e: out <= 12'h088;
      20'h0ad0f: out <= 12'h088;
      20'h0ad10: out <= 12'h088;
      20'h0ad11: out <= 12'h088;
      20'h0ad12: out <= 12'h088;
      20'h0ad13: out <= 12'h088;
      20'h0ad14: out <= 12'h088;
      20'h0ad15: out <= 12'h088;
      20'h0ad16: out <= 12'h088;
      20'h0ad17: out <= 12'h088;
      20'h0ad18: out <= 12'h088;
      20'h0ad19: out <= 12'h088;
      20'h0ad1a: out <= 12'h088;
      20'h0ad1b: out <= 12'h088;
      20'h0ad1c: out <= 12'h088;
      20'h0ad1d: out <= 12'h088;
      20'h0ad1e: out <= 12'h088;
      20'h0ad1f: out <= 12'h088;
      20'h0ad20: out <= 12'h088;
      20'h0ad21: out <= 12'h088;
      20'h0ad22: out <= 12'h088;
      20'h0ad23: out <= 12'h088;
      20'h0ad24: out <= 12'h088;
      20'h0ad25: out <= 12'h088;
      20'h0ad26: out <= 12'h088;
      20'h0ad27: out <= 12'h088;
      20'h0ad28: out <= 12'h088;
      20'h0ad29: out <= 12'h088;
      20'h0ad2a: out <= 12'h088;
      20'h0ad2b: out <= 12'h088;
      20'h0ad2c: out <= 12'h088;
      20'h0ad2d: out <= 12'h088;
      20'h0ad2e: out <= 12'h088;
      20'h0ad2f: out <= 12'h088;
      20'h0ad30: out <= 12'h088;
      20'h0ad31: out <= 12'h088;
      20'h0ad32: out <= 12'h088;
      20'h0ad33: out <= 12'h088;
      20'h0ad34: out <= 12'h088;
      20'h0ad35: out <= 12'h088;
      20'h0ad36: out <= 12'h088;
      20'h0ad37: out <= 12'h088;
      20'h0ad38: out <= 12'h088;
      20'h0ad39: out <= 12'hbb0;
      20'h0ad3a: out <= 12'h660;
      20'h0ad3b: out <= 12'h660;
      20'h0ad3c: out <= 12'h000;
      20'h0ad3d: out <= 12'hbb0;
      20'h0ad3e: out <= 12'hee9;
      20'h0ad3f: out <= 12'h660;
      20'h0ad40: out <= 12'h222;
      20'h0ad41: out <= 12'h660;
      20'h0ad42: out <= 12'hee9;
      20'h0ad43: out <= 12'hbb0;
      20'h0ad44: out <= 12'h222;
      20'h0ad45: out <= 12'hbb0;
      20'h0ad46: out <= 12'hee9;
      20'h0ad47: out <= 12'h660;
      20'h0ad48: out <= 12'hee9;
      20'h0ad49: out <= 12'hbb0;
      20'h0ad4a: out <= 12'h660;
      20'h0ad4b: out <= 12'h660;
      20'h0ad4c: out <= 12'h222;
      20'h0ad4d: out <= 12'hbb0;
      20'h0ad4e: out <= 12'h660;
      20'h0ad4f: out <= 12'h660;
      20'h0ad50: out <= 12'h603;
      20'h0ad51: out <= 12'h603;
      20'h0ad52: out <= 12'h603;
      20'h0ad53: out <= 12'h603;
      20'h0ad54: out <= 12'h000;
      20'h0ad55: out <= 12'hbbb;
      20'h0ad56: out <= 12'hbbb;
      20'h0ad57: out <= 12'hbbb;
      20'h0ad58: out <= 12'hbbb;
      20'h0ad59: out <= 12'hbbb;
      20'h0ad5a: out <= 12'h000;
      20'h0ad5b: out <= 12'h000;
      20'h0ad5c: out <= 12'h000;
      20'h0ad5d: out <= 12'h000;
      20'h0ad5e: out <= 12'h000;
      20'h0ad5f: out <= 12'hbbb;
      20'h0ad60: out <= 12'hbbb;
      20'h0ad61: out <= 12'h000;
      20'h0ad62: out <= 12'h000;
      20'h0ad63: out <= 12'h000;
      20'h0ad64: out <= 12'hbbb;
      20'h0ad65: out <= 12'hbbb;
      20'h0ad66: out <= 12'hbbb;
      20'h0ad67: out <= 12'hbbb;
      20'h0ad68: out <= 12'hbbb;
      20'h0ad69: out <= 12'hbbb;
      20'h0ad6a: out <= 12'hbbb;
      20'h0ad6b: out <= 12'h000;
      20'h0ad6c: out <= 12'h000;
      20'h0ad6d: out <= 12'hbbb;
      20'h0ad6e: out <= 12'hbbb;
      20'h0ad6f: out <= 12'hbbb;
      20'h0ad70: out <= 12'hbbb;
      20'h0ad71: out <= 12'hbbb;
      20'h0ad72: out <= 12'h000;
      20'h0ad73: out <= 12'h000;
      20'h0ad74: out <= 12'h000;
      20'h0ad75: out <= 12'h000;
      20'h0ad76: out <= 12'h000;
      20'h0ad77: out <= 12'h000;
      20'h0ad78: out <= 12'hbbb;
      20'h0ad79: out <= 12'hbbb;
      20'h0ad7a: out <= 12'h000;
      20'h0ad7b: out <= 12'h000;
      20'h0ad7c: out <= 12'h000;
      20'h0ad7d: out <= 12'hbbb;
      20'h0ad7e: out <= 12'hbbb;
      20'h0ad7f: out <= 12'hbbb;
      20'h0ad80: out <= 12'hbbb;
      20'h0ad81: out <= 12'hbbb;
      20'h0ad82: out <= 12'h000;
      20'h0ad83: out <= 12'h000;
      20'h0ad84: out <= 12'h000;
      20'h0ad85: out <= 12'hbbb;
      20'h0ad86: out <= 12'hbbb;
      20'h0ad87: out <= 12'hbbb;
      20'h0ad88: out <= 12'hbbb;
      20'h0ad89: out <= 12'hbbb;
      20'h0ad8a: out <= 12'h000;
      20'h0ad8b: out <= 12'h000;
      20'h0ad8c: out <= 12'h000;
      20'h0ad8d: out <= 12'h000;
      20'h0ad8e: out <= 12'hbbb;
      20'h0ad8f: out <= 12'hbbb;
      20'h0ad90: out <= 12'h000;
      20'h0ad91: out <= 12'h000;
      20'h0ad92: out <= 12'h000;
      20'h0ad93: out <= 12'h000;
      20'h0ad94: out <= 12'h000;
      20'h0ad95: out <= 12'hbbb;
      20'h0ad96: out <= 12'hbbb;
      20'h0ad97: out <= 12'hbbb;
      20'h0ad98: out <= 12'hbbb;
      20'h0ad99: out <= 12'hbbb;
      20'h0ad9a: out <= 12'h000;
      20'h0ad9b: out <= 12'h000;
      20'h0ad9c: out <= 12'h000;
      20'h0ad9d: out <= 12'hbbb;
      20'h0ad9e: out <= 12'hbbb;
      20'h0ad9f: out <= 12'hbbb;
      20'h0ada0: out <= 12'hbbb;
      20'h0ada1: out <= 12'h000;
      20'h0ada2: out <= 12'h000;
      20'h0ada3: out <= 12'h000;
      20'h0ada4: out <= 12'h603;
      20'h0ada5: out <= 12'h603;
      20'h0ada6: out <= 12'h603;
      20'h0ada7: out <= 12'h603;
      20'h0ada8: out <= 12'hee9;
      20'h0ada9: out <= 12'hf87;
      20'h0adaa: out <= 12'hf87;
      20'h0adab: out <= 12'hf87;
      20'h0adac: out <= 12'hf87;
      20'h0adad: out <= 12'hf87;
      20'h0adae: out <= 12'hf87;
      20'h0adaf: out <= 12'hb27;
      20'h0adb0: out <= 12'h000;
      20'h0adb1: out <= 12'h000;
      20'h0adb2: out <= 12'h000;
      20'h0adb3: out <= 12'h000;
      20'h0adb4: out <= 12'h000;
      20'h0adb5: out <= 12'h000;
      20'h0adb6: out <= 12'h000;
      20'h0adb7: out <= 12'h000;
      20'h0adb8: out <= 12'hfa9;
      20'h0adb9: out <= 12'hfa9;
      20'h0adba: out <= 12'hfa9;
      20'h0adbb: out <= 12'hfa9;
      20'h0adbc: out <= 12'hfa9;
      20'h0adbd: out <= 12'hfa9;
      20'h0adbe: out <= 12'hfa9;
      20'h0adbf: out <= 12'hfa9;
      20'h0adc0: out <= 12'hf76;
      20'h0adc1: out <= 12'hf76;
      20'h0adc2: out <= 12'hf76;
      20'h0adc3: out <= 12'hf76;
      20'h0adc4: out <= 12'hf76;
      20'h0adc5: out <= 12'hf76;
      20'h0adc6: out <= 12'hf76;
      20'h0adc7: out <= 12'hf76;
      20'h0adc8: out <= 12'hfa9;
      20'h0adc9: out <= 12'hfa9;
      20'h0adca: out <= 12'hfa9;
      20'h0adcb: out <= 12'hfa9;
      20'h0adcc: out <= 12'hfa9;
      20'h0adcd: out <= 12'hfa9;
      20'h0adce: out <= 12'hfa9;
      20'h0adcf: out <= 12'hfa9;
      20'h0add0: out <= 12'hf76;
      20'h0add1: out <= 12'hf76;
      20'h0add2: out <= 12'hf76;
      20'h0add3: out <= 12'hf76;
      20'h0add4: out <= 12'hf76;
      20'h0add5: out <= 12'hf76;
      20'h0add6: out <= 12'hf76;
      20'h0add7: out <= 12'hf76;
      20'h0add8: out <= 12'hfa9;
      20'h0add9: out <= 12'hfa9;
      20'h0adda: out <= 12'hfa9;
      20'h0addb: out <= 12'hfa9;
      20'h0addc: out <= 12'hfa9;
      20'h0addd: out <= 12'hfa9;
      20'h0adde: out <= 12'hfa9;
      20'h0addf: out <= 12'hfa9;
      20'h0ade0: out <= 12'h000;
      20'h0ade1: out <= 12'h000;
      20'h0ade2: out <= 12'h000;
      20'h0ade3: out <= 12'h000;
      20'h0ade4: out <= 12'h000;
      20'h0ade5: out <= 12'h000;
      20'h0ade6: out <= 12'h000;
      20'h0ade7: out <= 12'h000;
      20'h0ade8: out <= 12'h088;
      20'h0ade9: out <= 12'h088;
      20'h0adea: out <= 12'h088;
      20'h0adeb: out <= 12'h088;
      20'h0adec: out <= 12'h088;
      20'h0aded: out <= 12'h088;
      20'h0adee: out <= 12'h088;
      20'h0adef: out <= 12'h088;
      20'h0adf0: out <= 12'h088;
      20'h0adf1: out <= 12'h088;
      20'h0adf2: out <= 12'h088;
      20'h0adf3: out <= 12'h088;
      20'h0adf4: out <= 12'h088;
      20'h0adf5: out <= 12'h088;
      20'h0adf6: out <= 12'h088;
      20'h0adf7: out <= 12'h088;
      20'h0adf8: out <= 12'h088;
      20'h0adf9: out <= 12'h088;
      20'h0adfa: out <= 12'h088;
      20'h0adfb: out <= 12'h088;
      20'h0adfc: out <= 12'h088;
      20'h0adfd: out <= 12'h088;
      20'h0adfe: out <= 12'h088;
      20'h0adff: out <= 12'h088;
      20'h0ae00: out <= 12'h088;
      20'h0ae01: out <= 12'h088;
      20'h0ae02: out <= 12'h088;
      20'h0ae03: out <= 12'h088;
      20'h0ae04: out <= 12'h088;
      20'h0ae05: out <= 12'h088;
      20'h0ae06: out <= 12'h088;
      20'h0ae07: out <= 12'h088;
      20'h0ae08: out <= 12'h088;
      20'h0ae09: out <= 12'h088;
      20'h0ae0a: out <= 12'h088;
      20'h0ae0b: out <= 12'h088;
      20'h0ae0c: out <= 12'h088;
      20'h0ae0d: out <= 12'h088;
      20'h0ae0e: out <= 12'h088;
      20'h0ae0f: out <= 12'h088;
      20'h0ae10: out <= 12'h088;
      20'h0ae11: out <= 12'h088;
      20'h0ae12: out <= 12'h088;
      20'h0ae13: out <= 12'h088;
      20'h0ae14: out <= 12'h088;
      20'h0ae15: out <= 12'h088;
      20'h0ae16: out <= 12'h088;
      20'h0ae17: out <= 12'h088;
      20'h0ae18: out <= 12'h088;
      20'h0ae19: out <= 12'h088;
      20'h0ae1a: out <= 12'h088;
      20'h0ae1b: out <= 12'h088;
      20'h0ae1c: out <= 12'h088;
      20'h0ae1d: out <= 12'h088;
      20'h0ae1e: out <= 12'h088;
      20'h0ae1f: out <= 12'h088;
      20'h0ae20: out <= 12'h088;
      20'h0ae21: out <= 12'h088;
      20'h0ae22: out <= 12'h088;
      20'h0ae23: out <= 12'h088;
      20'h0ae24: out <= 12'h088;
      20'h0ae25: out <= 12'h088;
      20'h0ae26: out <= 12'h088;
      20'h0ae27: out <= 12'h088;
      20'h0ae28: out <= 12'h088;
      20'h0ae29: out <= 12'h088;
      20'h0ae2a: out <= 12'h088;
      20'h0ae2b: out <= 12'h088;
      20'h0ae2c: out <= 12'h088;
      20'h0ae2d: out <= 12'h088;
      20'h0ae2e: out <= 12'h088;
      20'h0ae2f: out <= 12'h088;
      20'h0ae30: out <= 12'h088;
      20'h0ae31: out <= 12'h088;
      20'h0ae32: out <= 12'h088;
      20'h0ae33: out <= 12'h088;
      20'h0ae34: out <= 12'h088;
      20'h0ae35: out <= 12'h088;
      20'h0ae36: out <= 12'h088;
      20'h0ae37: out <= 12'h088;
      20'h0ae38: out <= 12'h088;
      20'h0ae39: out <= 12'h088;
      20'h0ae3a: out <= 12'h088;
      20'h0ae3b: out <= 12'h088;
      20'h0ae3c: out <= 12'h088;
      20'h0ae3d: out <= 12'h088;
      20'h0ae3e: out <= 12'h088;
      20'h0ae3f: out <= 12'h088;
      20'h0ae40: out <= 12'h088;
      20'h0ae41: out <= 12'h088;
      20'h0ae42: out <= 12'h088;
      20'h0ae43: out <= 12'h088;
      20'h0ae44: out <= 12'h088;
      20'h0ae45: out <= 12'h088;
      20'h0ae46: out <= 12'h088;
      20'h0ae47: out <= 12'h088;
      20'h0ae48: out <= 12'h088;
      20'h0ae49: out <= 12'h088;
      20'h0ae4a: out <= 12'h088;
      20'h0ae4b: out <= 12'h088;
      20'h0ae4c: out <= 12'h088;
      20'h0ae4d: out <= 12'h088;
      20'h0ae4e: out <= 12'h088;
      20'h0ae4f: out <= 12'h088;
      20'h0ae50: out <= 12'h088;
      20'h0ae51: out <= 12'hbb0;
      20'h0ae52: out <= 12'h000;
      20'h0ae53: out <= 12'h000;
      20'h0ae54: out <= 12'h000;
      20'h0ae55: out <= 12'h000;
      20'h0ae56: out <= 12'h000;
      20'h0ae57: out <= 12'h000;
      20'h0ae58: out <= 12'h222;
      20'h0ae59: out <= 12'h222;
      20'h0ae5a: out <= 12'h222;
      20'h0ae5b: out <= 12'h222;
      20'h0ae5c: out <= 12'h222;
      20'h0ae5d: out <= 12'h222;
      20'h0ae5e: out <= 12'h222;
      20'h0ae5f: out <= 12'h660;
      20'h0ae60: out <= 12'hee9;
      20'h0ae61: out <= 12'hbb0;
      20'h0ae62: out <= 12'h222;
      20'h0ae63: out <= 12'h222;
      20'h0ae64: out <= 12'h222;
      20'h0ae65: out <= 12'h222;
      20'h0ae66: out <= 12'h222;
      20'h0ae67: out <= 12'h222;
      20'h0ae68: out <= 12'h603;
      20'h0ae69: out <= 12'h603;
      20'h0ae6a: out <= 12'h603;
      20'h0ae6b: out <= 12'h603;
      20'h0ae6c: out <= 12'h000;
      20'h0ae6d: out <= 12'h000;
      20'h0ae6e: out <= 12'h000;
      20'h0ae6f: out <= 12'h000;
      20'h0ae70: out <= 12'h000;
      20'h0ae71: out <= 12'h000;
      20'h0ae72: out <= 12'h000;
      20'h0ae73: out <= 12'h000;
      20'h0ae74: out <= 12'h000;
      20'h0ae75: out <= 12'h000;
      20'h0ae76: out <= 12'h000;
      20'h0ae77: out <= 12'h000;
      20'h0ae78: out <= 12'h000;
      20'h0ae79: out <= 12'h000;
      20'h0ae7a: out <= 12'h000;
      20'h0ae7b: out <= 12'h000;
      20'h0ae7c: out <= 12'h000;
      20'h0ae7d: out <= 12'h000;
      20'h0ae7e: out <= 12'h000;
      20'h0ae7f: out <= 12'h000;
      20'h0ae80: out <= 12'h000;
      20'h0ae81: out <= 12'h000;
      20'h0ae82: out <= 12'h000;
      20'h0ae83: out <= 12'h000;
      20'h0ae84: out <= 12'h000;
      20'h0ae85: out <= 12'h000;
      20'h0ae86: out <= 12'h000;
      20'h0ae87: out <= 12'h000;
      20'h0ae88: out <= 12'h000;
      20'h0ae89: out <= 12'h000;
      20'h0ae8a: out <= 12'h000;
      20'h0ae8b: out <= 12'h000;
      20'h0ae8c: out <= 12'h000;
      20'h0ae8d: out <= 12'h000;
      20'h0ae8e: out <= 12'h000;
      20'h0ae8f: out <= 12'h000;
      20'h0ae90: out <= 12'h000;
      20'h0ae91: out <= 12'h000;
      20'h0ae92: out <= 12'h000;
      20'h0ae93: out <= 12'h000;
      20'h0ae94: out <= 12'h000;
      20'h0ae95: out <= 12'h000;
      20'h0ae96: out <= 12'h000;
      20'h0ae97: out <= 12'h000;
      20'h0ae98: out <= 12'h000;
      20'h0ae99: out <= 12'h000;
      20'h0ae9a: out <= 12'h000;
      20'h0ae9b: out <= 12'h000;
      20'h0ae9c: out <= 12'h000;
      20'h0ae9d: out <= 12'h000;
      20'h0ae9e: out <= 12'h000;
      20'h0ae9f: out <= 12'h000;
      20'h0aea0: out <= 12'h000;
      20'h0aea1: out <= 12'h000;
      20'h0aea2: out <= 12'h000;
      20'h0aea3: out <= 12'h000;
      20'h0aea4: out <= 12'h000;
      20'h0aea5: out <= 12'h000;
      20'h0aea6: out <= 12'h000;
      20'h0aea7: out <= 12'h000;
      20'h0aea8: out <= 12'h000;
      20'h0aea9: out <= 12'h000;
      20'h0aeaa: out <= 12'h000;
      20'h0aeab: out <= 12'h000;
      20'h0aeac: out <= 12'h000;
      20'h0aead: out <= 12'h000;
      20'h0aeae: out <= 12'h000;
      20'h0aeaf: out <= 12'h000;
      20'h0aeb0: out <= 12'h000;
      20'h0aeb1: out <= 12'h000;
      20'h0aeb2: out <= 12'h000;
      20'h0aeb3: out <= 12'h000;
      20'h0aeb4: out <= 12'h000;
      20'h0aeb5: out <= 12'h000;
      20'h0aeb6: out <= 12'h000;
      20'h0aeb7: out <= 12'h000;
      20'h0aeb8: out <= 12'h000;
      20'h0aeb9: out <= 12'h000;
      20'h0aeba: out <= 12'h000;
      20'h0aebb: out <= 12'h000;
      20'h0aebc: out <= 12'h603;
      20'h0aebd: out <= 12'h603;
      20'h0aebe: out <= 12'h603;
      20'h0aebf: out <= 12'h603;
      20'h0aec0: out <= 12'hb27;
      20'h0aec1: out <= 12'hb27;
      20'h0aec2: out <= 12'hb27;
      20'h0aec3: out <= 12'hb27;
      20'h0aec4: out <= 12'hb27;
      20'h0aec5: out <= 12'hb27;
      20'h0aec6: out <= 12'hb27;
      20'h0aec7: out <= 12'hb27;
      20'h0aec8: out <= 12'h000;
      20'h0aec9: out <= 12'h000;
      20'h0aeca: out <= 12'h000;
      20'h0aecb: out <= 12'h000;
      20'h0aecc: out <= 12'h000;
      20'h0aecd: out <= 12'h000;
      20'h0aece: out <= 12'h000;
      20'h0aecf: out <= 12'h000;
      20'h0aed0: out <= 12'hfa9;
      20'h0aed1: out <= 12'hfa9;
      20'h0aed2: out <= 12'hfa9;
      20'h0aed3: out <= 12'hfa9;
      20'h0aed4: out <= 12'hfa9;
      20'h0aed5: out <= 12'hfa9;
      20'h0aed6: out <= 12'hfa9;
      20'h0aed7: out <= 12'hfa9;
      20'h0aed8: out <= 12'hf76;
      20'h0aed9: out <= 12'hf76;
      20'h0aeda: out <= 12'hf76;
      20'h0aedb: out <= 12'hf76;
      20'h0aedc: out <= 12'hf76;
      20'h0aedd: out <= 12'hf76;
      20'h0aede: out <= 12'hf76;
      20'h0aedf: out <= 12'hf76;
      20'h0aee0: out <= 12'hfa9;
      20'h0aee1: out <= 12'hfa9;
      20'h0aee2: out <= 12'hfa9;
      20'h0aee3: out <= 12'hfa9;
      20'h0aee4: out <= 12'hfa9;
      20'h0aee5: out <= 12'hfa9;
      20'h0aee6: out <= 12'hfa9;
      20'h0aee7: out <= 12'hfa9;
      20'h0aee8: out <= 12'hf76;
      20'h0aee9: out <= 12'hf76;
      20'h0aeea: out <= 12'hf76;
      20'h0aeeb: out <= 12'hf76;
      20'h0aeec: out <= 12'hf76;
      20'h0aeed: out <= 12'hf76;
      20'h0aeee: out <= 12'hf76;
      20'h0aeef: out <= 12'hf76;
      20'h0aef0: out <= 12'hfa9;
      20'h0aef1: out <= 12'hfa9;
      20'h0aef2: out <= 12'hfa9;
      20'h0aef3: out <= 12'hfa9;
      20'h0aef4: out <= 12'hfa9;
      20'h0aef5: out <= 12'hfa9;
      20'h0aef6: out <= 12'hfa9;
      20'h0aef7: out <= 12'hfa9;
      20'h0aef8: out <= 12'h000;
      20'h0aef9: out <= 12'h000;
      20'h0aefa: out <= 12'h000;
      20'h0aefb: out <= 12'h000;
      20'h0aefc: out <= 12'h000;
      20'h0aefd: out <= 12'h000;
      20'h0aefe: out <= 12'h000;
      20'h0aeff: out <= 12'h000;
      20'h0af00: out <= 12'h088;
      20'h0af01: out <= 12'h088;
      20'h0af02: out <= 12'h088;
      20'h0af03: out <= 12'h088;
      20'h0af04: out <= 12'h088;
      20'h0af05: out <= 12'h088;
      20'h0af06: out <= 12'h088;
      20'h0af07: out <= 12'h088;
      20'h0af08: out <= 12'h088;
      20'h0af09: out <= 12'h088;
      20'h0af0a: out <= 12'h088;
      20'h0af0b: out <= 12'h088;
      20'h0af0c: out <= 12'h088;
      20'h0af0d: out <= 12'h088;
      20'h0af0e: out <= 12'h088;
      20'h0af0f: out <= 12'h088;
      20'h0af10: out <= 12'h088;
      20'h0af11: out <= 12'h088;
      20'h0af12: out <= 12'h088;
      20'h0af13: out <= 12'h088;
      20'h0af14: out <= 12'h088;
      20'h0af15: out <= 12'h088;
      20'h0af16: out <= 12'h088;
      20'h0af17: out <= 12'h088;
      20'h0af18: out <= 12'h088;
      20'h0af19: out <= 12'h088;
      20'h0af1a: out <= 12'h088;
      20'h0af1b: out <= 12'h088;
      20'h0af1c: out <= 12'h088;
      20'h0af1d: out <= 12'h088;
      20'h0af1e: out <= 12'h088;
      20'h0af1f: out <= 12'h088;
      20'h0af20: out <= 12'h088;
      20'h0af21: out <= 12'h088;
      20'h0af22: out <= 12'h088;
      20'h0af23: out <= 12'h088;
      20'h0af24: out <= 12'h088;
      20'h0af25: out <= 12'h088;
      20'h0af26: out <= 12'h088;
      20'h0af27: out <= 12'h088;
      20'h0af28: out <= 12'h088;
      20'h0af29: out <= 12'h088;
      20'h0af2a: out <= 12'h088;
      20'h0af2b: out <= 12'h088;
      20'h0af2c: out <= 12'h088;
      20'h0af2d: out <= 12'h088;
      20'h0af2e: out <= 12'h088;
      20'h0af2f: out <= 12'h088;
      20'h0af30: out <= 12'h088;
      20'h0af31: out <= 12'h088;
      20'h0af32: out <= 12'h088;
      20'h0af33: out <= 12'h088;
      20'h0af34: out <= 12'h088;
      20'h0af35: out <= 12'h088;
      20'h0af36: out <= 12'h088;
      20'h0af37: out <= 12'h088;
      20'h0af38: out <= 12'h088;
      20'h0af39: out <= 12'h088;
      20'h0af3a: out <= 12'h088;
      20'h0af3b: out <= 12'h088;
      20'h0af3c: out <= 12'h088;
      20'h0af3d: out <= 12'h088;
      20'h0af3e: out <= 12'h088;
      20'h0af3f: out <= 12'h088;
      20'h0af40: out <= 12'h088;
      20'h0af41: out <= 12'h088;
      20'h0af42: out <= 12'h088;
      20'h0af43: out <= 12'h088;
      20'h0af44: out <= 12'h088;
      20'h0af45: out <= 12'h088;
      20'h0af46: out <= 12'h088;
      20'h0af47: out <= 12'h088;
      20'h0af48: out <= 12'h088;
      20'h0af49: out <= 12'h088;
      20'h0af4a: out <= 12'h088;
      20'h0af4b: out <= 12'h088;
      20'h0af4c: out <= 12'h088;
      20'h0af4d: out <= 12'h088;
      20'h0af4e: out <= 12'h088;
      20'h0af4f: out <= 12'h088;
      20'h0af50: out <= 12'h088;
      20'h0af51: out <= 12'h088;
      20'h0af52: out <= 12'h088;
      20'h0af53: out <= 12'h088;
      20'h0af54: out <= 12'h088;
      20'h0af55: out <= 12'h088;
      20'h0af56: out <= 12'h088;
      20'h0af57: out <= 12'h088;
      20'h0af58: out <= 12'h088;
      20'h0af59: out <= 12'h088;
      20'h0af5a: out <= 12'h088;
      20'h0af5b: out <= 12'h088;
      20'h0af5c: out <= 12'h088;
      20'h0af5d: out <= 12'h088;
      20'h0af5e: out <= 12'h088;
      20'h0af5f: out <= 12'h088;
      20'h0af60: out <= 12'h088;
      20'h0af61: out <= 12'h088;
      20'h0af62: out <= 12'h088;
      20'h0af63: out <= 12'h088;
      20'h0af64: out <= 12'h088;
      20'h0af65: out <= 12'h088;
      20'h0af66: out <= 12'h088;
      20'h0af67: out <= 12'h088;
      20'h0af68: out <= 12'h088;
      20'h0af69: out <= 12'h603;
      20'h0af6a: out <= 12'h603;
      20'h0af6b: out <= 12'h603;
      20'h0af6c: out <= 12'h603;
      20'h0af6d: out <= 12'h603;
      20'h0af6e: out <= 12'h603;
      20'h0af6f: out <= 12'h603;
      20'h0af70: out <= 12'h603;
      20'h0af71: out <= 12'h603;
      20'h0af72: out <= 12'h603;
      20'h0af73: out <= 12'h603;
      20'h0af74: out <= 12'h603;
      20'h0af75: out <= 12'h603;
      20'h0af76: out <= 12'h603;
      20'h0af77: out <= 12'h603;
      20'h0af78: out <= 12'h603;
      20'h0af79: out <= 12'h603;
      20'h0af7a: out <= 12'h603;
      20'h0af7b: out <= 12'h603;
      20'h0af7c: out <= 12'h603;
      20'h0af7d: out <= 12'h603;
      20'h0af7e: out <= 12'h603;
      20'h0af7f: out <= 12'h603;
      20'h0af80: out <= 12'h603;
      20'h0af81: out <= 12'h603;
      20'h0af82: out <= 12'h603;
      20'h0af83: out <= 12'h603;
      20'h0af84: out <= 12'h000;
      20'h0af85: out <= 12'h8d0;
      20'h0af86: out <= 12'h8d0;
      20'h0af87: out <= 12'h8d0;
      20'h0af88: out <= 12'h8d0;
      20'h0af89: out <= 12'h8d0;
      20'h0af8a: out <= 12'h000;
      20'h0af8b: out <= 12'h000;
      20'h0af8c: out <= 12'h000;
      20'h0af8d: out <= 12'h000;
      20'h0af8e: out <= 12'h000;
      20'h0af8f: out <= 12'h8d0;
      20'h0af90: out <= 12'h8d0;
      20'h0af91: out <= 12'h000;
      20'h0af92: out <= 12'h000;
      20'h0af93: out <= 12'h000;
      20'h0af94: out <= 12'h000;
      20'h0af95: out <= 12'h8d0;
      20'h0af96: out <= 12'h8d0;
      20'h0af97: out <= 12'h8d0;
      20'h0af98: out <= 12'h8d0;
      20'h0af99: out <= 12'h8d0;
      20'h0af9a: out <= 12'h000;
      20'h0af9b: out <= 12'h000;
      20'h0af9c: out <= 12'h000;
      20'h0af9d: out <= 12'h8d0;
      20'h0af9e: out <= 12'h8d0;
      20'h0af9f: out <= 12'h8d0;
      20'h0afa0: out <= 12'h8d0;
      20'h0afa1: out <= 12'h8d0;
      20'h0afa2: out <= 12'h000;
      20'h0afa3: out <= 12'h000;
      20'h0afa4: out <= 12'h000;
      20'h0afa5: out <= 12'h000;
      20'h0afa6: out <= 12'h000;
      20'h0afa7: out <= 12'h8d0;
      20'h0afa8: out <= 12'h8d0;
      20'h0afa9: out <= 12'h8d0;
      20'h0afaa: out <= 12'h000;
      20'h0afab: out <= 12'h000;
      20'h0afac: out <= 12'h8d0;
      20'h0afad: out <= 12'h8d0;
      20'h0afae: out <= 12'h8d0;
      20'h0afaf: out <= 12'h8d0;
      20'h0afb0: out <= 12'h8d0;
      20'h0afb1: out <= 12'h8d0;
      20'h0afb2: out <= 12'h8d0;
      20'h0afb3: out <= 12'h000;
      20'h0afb4: out <= 12'h000;
      20'h0afb5: out <= 12'h000;
      20'h0afb6: out <= 12'h8d0;
      20'h0afb7: out <= 12'h8d0;
      20'h0afb8: out <= 12'h8d0;
      20'h0afb9: out <= 12'h8d0;
      20'h0afba: out <= 12'h000;
      20'h0afbb: out <= 12'h000;
      20'h0afbc: out <= 12'h8d0;
      20'h0afbd: out <= 12'h8d0;
      20'h0afbe: out <= 12'h8d0;
      20'h0afbf: out <= 12'h8d0;
      20'h0afc0: out <= 12'h8d0;
      20'h0afc1: out <= 12'h8d0;
      20'h0afc2: out <= 12'h8d0;
      20'h0afc3: out <= 12'h000;
      20'h0afc4: out <= 12'h000;
      20'h0afc5: out <= 12'h8d0;
      20'h0afc6: out <= 12'h8d0;
      20'h0afc7: out <= 12'h8d0;
      20'h0afc8: out <= 12'h8d0;
      20'h0afc9: out <= 12'h8d0;
      20'h0afca: out <= 12'h000;
      20'h0afcb: out <= 12'h000;
      20'h0afcc: out <= 12'h000;
      20'h0afcd: out <= 12'h8d0;
      20'h0afce: out <= 12'h8d0;
      20'h0afcf: out <= 12'h8d0;
      20'h0afd0: out <= 12'h8d0;
      20'h0afd1: out <= 12'h8d0;
      20'h0afd2: out <= 12'h000;
      20'h0afd3: out <= 12'h000;
      20'h0afd4: out <= 12'h603;
      20'h0afd5: out <= 12'h603;
      20'h0afd6: out <= 12'h603;
      20'h0afd7: out <= 12'h603;
      20'h0afd8: out <= 12'hee9;
      20'h0afd9: out <= 12'hee9;
      20'h0afda: out <= 12'hee9;
      20'h0afdb: out <= 12'hee9;
      20'h0afdc: out <= 12'hee9;
      20'h0afdd: out <= 12'hee9;
      20'h0afde: out <= 12'hee9;
      20'h0afdf: out <= 12'hb27;
      20'h0afe0: out <= 12'h000;
      20'h0afe1: out <= 12'h000;
      20'h0afe2: out <= 12'h000;
      20'h0afe3: out <= 12'h000;
      20'h0afe4: out <= 12'h000;
      20'h0afe5: out <= 12'h000;
      20'h0afe6: out <= 12'h000;
      20'h0afe7: out <= 12'h000;
      20'h0afe8: out <= 12'h777;
      20'h0afe9: out <= 12'h777;
      20'h0afea: out <= 12'h777;
      20'h0afeb: out <= 12'h777;
      20'h0afec: out <= 12'h777;
      20'h0afed: out <= 12'h777;
      20'h0afee: out <= 12'h777;
      20'h0afef: out <= 12'h777;
      20'h0aff0: out <= 12'h777;
      20'h0aff1: out <= 12'h777;
      20'h0aff2: out <= 12'h777;
      20'h0aff3: out <= 12'h777;
      20'h0aff4: out <= 12'h777;
      20'h0aff5: out <= 12'h777;
      20'h0aff6: out <= 12'h777;
      20'h0aff7: out <= 12'h777;
      20'h0aff8: out <= 12'h000;
      20'h0aff9: out <= 12'h000;
      20'h0affa: out <= 12'h000;
      20'h0affb: out <= 12'h000;
      20'h0affc: out <= 12'h000;
      20'h0affd: out <= 12'h000;
      20'h0affe: out <= 12'h000;
      20'h0afff: out <= 12'h000;
      20'h0b000: out <= 12'h000;
      20'h0b001: out <= 12'h000;
      20'h0b002: out <= 12'h000;
      20'h0b003: out <= 12'h000;
      20'h0b004: out <= 12'h000;
      20'h0b005: out <= 12'h000;
      20'h0b006: out <= 12'h000;
      20'h0b007: out <= 12'h000;
      20'h0b008: out <= 12'h000;
      20'h0b009: out <= 12'h000;
      20'h0b00a: out <= 12'h000;
      20'h0b00b: out <= 12'h000;
      20'h0b00c: out <= 12'h000;
      20'h0b00d: out <= 12'h000;
      20'h0b00e: out <= 12'h000;
      20'h0b00f: out <= 12'h000;
      20'h0b010: out <= 12'h000;
      20'h0b011: out <= 12'h000;
      20'h0b012: out <= 12'h000;
      20'h0b013: out <= 12'h000;
      20'h0b014: out <= 12'h000;
      20'h0b015: out <= 12'h000;
      20'h0b016: out <= 12'h000;
      20'h0b017: out <= 12'h000;
      20'h0b018: out <= 12'h088;
      20'h0b019: out <= 12'h088;
      20'h0b01a: out <= 12'h088;
      20'h0b01b: out <= 12'h088;
      20'h0b01c: out <= 12'h088;
      20'h0b01d: out <= 12'h088;
      20'h0b01e: out <= 12'h088;
      20'h0b01f: out <= 12'h088;
      20'h0b020: out <= 12'h088;
      20'h0b021: out <= 12'h088;
      20'h0b022: out <= 12'h088;
      20'h0b023: out <= 12'h088;
      20'h0b024: out <= 12'h088;
      20'h0b025: out <= 12'h088;
      20'h0b026: out <= 12'h088;
      20'h0b027: out <= 12'h088;
      20'h0b028: out <= 12'h088;
      20'h0b029: out <= 12'h088;
      20'h0b02a: out <= 12'h088;
      20'h0b02b: out <= 12'h088;
      20'h0b02c: out <= 12'h088;
      20'h0b02d: out <= 12'h088;
      20'h0b02e: out <= 12'h088;
      20'h0b02f: out <= 12'h088;
      20'h0b030: out <= 12'h088;
      20'h0b031: out <= 12'h088;
      20'h0b032: out <= 12'h088;
      20'h0b033: out <= 12'h088;
      20'h0b034: out <= 12'h088;
      20'h0b035: out <= 12'h088;
      20'h0b036: out <= 12'h088;
      20'h0b037: out <= 12'h088;
      20'h0b038: out <= 12'h088;
      20'h0b039: out <= 12'h088;
      20'h0b03a: out <= 12'h088;
      20'h0b03b: out <= 12'h088;
      20'h0b03c: out <= 12'h088;
      20'h0b03d: out <= 12'h088;
      20'h0b03e: out <= 12'h088;
      20'h0b03f: out <= 12'h088;
      20'h0b040: out <= 12'h088;
      20'h0b041: out <= 12'h088;
      20'h0b042: out <= 12'h088;
      20'h0b043: out <= 12'h088;
      20'h0b044: out <= 12'h088;
      20'h0b045: out <= 12'h088;
      20'h0b046: out <= 12'h088;
      20'h0b047: out <= 12'h088;
      20'h0b048: out <= 12'h088;
      20'h0b049: out <= 12'h088;
      20'h0b04a: out <= 12'h088;
      20'h0b04b: out <= 12'h088;
      20'h0b04c: out <= 12'h088;
      20'h0b04d: out <= 12'h088;
      20'h0b04e: out <= 12'h088;
      20'h0b04f: out <= 12'h088;
      20'h0b050: out <= 12'h088;
      20'h0b051: out <= 12'h088;
      20'h0b052: out <= 12'h088;
      20'h0b053: out <= 12'h088;
      20'h0b054: out <= 12'h088;
      20'h0b055: out <= 12'h088;
      20'h0b056: out <= 12'h088;
      20'h0b057: out <= 12'h088;
      20'h0b058: out <= 12'h088;
      20'h0b059: out <= 12'h088;
      20'h0b05a: out <= 12'h088;
      20'h0b05b: out <= 12'h088;
      20'h0b05c: out <= 12'h088;
      20'h0b05d: out <= 12'h088;
      20'h0b05e: out <= 12'h088;
      20'h0b05f: out <= 12'h088;
      20'h0b060: out <= 12'h088;
      20'h0b061: out <= 12'h088;
      20'h0b062: out <= 12'h088;
      20'h0b063: out <= 12'h088;
      20'h0b064: out <= 12'h088;
      20'h0b065: out <= 12'h088;
      20'h0b066: out <= 12'h088;
      20'h0b067: out <= 12'h088;
      20'h0b068: out <= 12'h088;
      20'h0b069: out <= 12'h088;
      20'h0b06a: out <= 12'h088;
      20'h0b06b: out <= 12'h088;
      20'h0b06c: out <= 12'h088;
      20'h0b06d: out <= 12'h088;
      20'h0b06e: out <= 12'h088;
      20'h0b06f: out <= 12'h088;
      20'h0b070: out <= 12'h088;
      20'h0b071: out <= 12'h088;
      20'h0b072: out <= 12'h088;
      20'h0b073: out <= 12'h088;
      20'h0b074: out <= 12'h088;
      20'h0b075: out <= 12'h088;
      20'h0b076: out <= 12'h088;
      20'h0b077: out <= 12'h088;
      20'h0b078: out <= 12'h088;
      20'h0b079: out <= 12'h088;
      20'h0b07a: out <= 12'h088;
      20'h0b07b: out <= 12'h088;
      20'h0b07c: out <= 12'h088;
      20'h0b07d: out <= 12'h088;
      20'h0b07e: out <= 12'h088;
      20'h0b07f: out <= 12'h088;
      20'h0b080: out <= 12'h088;
      20'h0b081: out <= 12'h603;
      20'h0b082: out <= 12'h603;
      20'h0b083: out <= 12'h603;
      20'h0b084: out <= 12'h603;
      20'h0b085: out <= 12'h603;
      20'h0b086: out <= 12'h603;
      20'h0b087: out <= 12'h603;
      20'h0b088: out <= 12'h603;
      20'h0b089: out <= 12'h603;
      20'h0b08a: out <= 12'h603;
      20'h0b08b: out <= 12'h603;
      20'h0b08c: out <= 12'h603;
      20'h0b08d: out <= 12'h603;
      20'h0b08e: out <= 12'h603;
      20'h0b08f: out <= 12'h603;
      20'h0b090: out <= 12'h603;
      20'h0b091: out <= 12'h603;
      20'h0b092: out <= 12'h603;
      20'h0b093: out <= 12'h603;
      20'h0b094: out <= 12'h603;
      20'h0b095: out <= 12'h603;
      20'h0b096: out <= 12'h603;
      20'h0b097: out <= 12'h603;
      20'h0b098: out <= 12'h603;
      20'h0b099: out <= 12'h603;
      20'h0b09a: out <= 12'h603;
      20'h0b09b: out <= 12'h603;
      20'h0b09c: out <= 12'h8d0;
      20'h0b09d: out <= 12'h8d0;
      20'h0b09e: out <= 12'h000;
      20'h0b09f: out <= 12'h000;
      20'h0b0a0: out <= 12'h000;
      20'h0b0a1: out <= 12'h8d0;
      20'h0b0a2: out <= 12'h8d0;
      20'h0b0a3: out <= 12'h000;
      20'h0b0a4: out <= 12'h000;
      20'h0b0a5: out <= 12'h000;
      20'h0b0a6: out <= 12'h8d0;
      20'h0b0a7: out <= 12'h8d0;
      20'h0b0a8: out <= 12'h8d0;
      20'h0b0a9: out <= 12'h000;
      20'h0b0aa: out <= 12'h000;
      20'h0b0ab: out <= 12'h000;
      20'h0b0ac: out <= 12'h8d0;
      20'h0b0ad: out <= 12'h8d0;
      20'h0b0ae: out <= 12'h000;
      20'h0b0af: out <= 12'h000;
      20'h0b0b0: out <= 12'h000;
      20'h0b0b1: out <= 12'h8d0;
      20'h0b0b2: out <= 12'h8d0;
      20'h0b0b3: out <= 12'h000;
      20'h0b0b4: out <= 12'h8d0;
      20'h0b0b5: out <= 12'h8d0;
      20'h0b0b6: out <= 12'h000;
      20'h0b0b7: out <= 12'h000;
      20'h0b0b8: out <= 12'h000;
      20'h0b0b9: out <= 12'h8d0;
      20'h0b0ba: out <= 12'h8d0;
      20'h0b0bb: out <= 12'h000;
      20'h0b0bc: out <= 12'h000;
      20'h0b0bd: out <= 12'h000;
      20'h0b0be: out <= 12'h8d0;
      20'h0b0bf: out <= 12'h8d0;
      20'h0b0c0: out <= 12'h8d0;
      20'h0b0c1: out <= 12'h8d0;
      20'h0b0c2: out <= 12'h000;
      20'h0b0c3: out <= 12'h000;
      20'h0b0c4: out <= 12'h8d0;
      20'h0b0c5: out <= 12'h8d0;
      20'h0b0c6: out <= 12'h000;
      20'h0b0c7: out <= 12'h000;
      20'h0b0c8: out <= 12'h000;
      20'h0b0c9: out <= 12'h000;
      20'h0b0ca: out <= 12'h000;
      20'h0b0cb: out <= 12'h000;
      20'h0b0cc: out <= 12'h000;
      20'h0b0cd: out <= 12'h8d0;
      20'h0b0ce: out <= 12'h8d0;
      20'h0b0cf: out <= 12'h000;
      20'h0b0d0: out <= 12'h000;
      20'h0b0d1: out <= 12'h000;
      20'h0b0d2: out <= 12'h000;
      20'h0b0d3: out <= 12'h000;
      20'h0b0d4: out <= 12'h8d0;
      20'h0b0d5: out <= 12'h8d0;
      20'h0b0d6: out <= 12'h000;
      20'h0b0d7: out <= 12'h000;
      20'h0b0d8: out <= 12'h000;
      20'h0b0d9: out <= 12'h8d0;
      20'h0b0da: out <= 12'h8d0;
      20'h0b0db: out <= 12'h000;
      20'h0b0dc: out <= 12'h8d0;
      20'h0b0dd: out <= 12'h8d0;
      20'h0b0de: out <= 12'h000;
      20'h0b0df: out <= 12'h000;
      20'h0b0e0: out <= 12'h000;
      20'h0b0e1: out <= 12'h8d0;
      20'h0b0e2: out <= 12'h8d0;
      20'h0b0e3: out <= 12'h000;
      20'h0b0e4: out <= 12'h8d0;
      20'h0b0e5: out <= 12'h8d0;
      20'h0b0e6: out <= 12'h000;
      20'h0b0e7: out <= 12'h000;
      20'h0b0e8: out <= 12'h000;
      20'h0b0e9: out <= 12'h8d0;
      20'h0b0ea: out <= 12'h8d0;
      20'h0b0eb: out <= 12'h000;
      20'h0b0ec: out <= 12'h603;
      20'h0b0ed: out <= 12'h603;
      20'h0b0ee: out <= 12'h603;
      20'h0b0ef: out <= 12'h603;
      20'h0b0f0: out <= 12'hee9;
      20'h0b0f1: out <= 12'hf87;
      20'h0b0f2: out <= 12'hf87;
      20'h0b0f3: out <= 12'hf87;
      20'h0b0f4: out <= 12'hf87;
      20'h0b0f5: out <= 12'hf87;
      20'h0b0f6: out <= 12'hf87;
      20'h0b0f7: out <= 12'hb27;
      20'h0b0f8: out <= 12'h000;
      20'h0b0f9: out <= 12'h000;
      20'h0b0fa: out <= 12'h000;
      20'h0b0fb: out <= 12'h000;
      20'h0b0fc: out <= 12'h000;
      20'h0b0fd: out <= 12'h000;
      20'h0b0fe: out <= 12'h000;
      20'h0b0ff: out <= 12'h000;
      20'h0b100: out <= 12'h777;
      20'h0b101: out <= 12'h777;
      20'h0b102: out <= 12'h555;
      20'h0b103: out <= 12'h555;
      20'h0b104: out <= 12'h555;
      20'h0b105: out <= 12'h555;
      20'h0b106: out <= 12'h555;
      20'h0b107: out <= 12'h555;
      20'h0b108: out <= 12'h555;
      20'h0b109: out <= 12'h555;
      20'h0b10a: out <= 12'h555;
      20'h0b10b: out <= 12'h555;
      20'h0b10c: out <= 12'h555;
      20'h0b10d: out <= 12'h555;
      20'h0b10e: out <= 12'h777;
      20'h0b10f: out <= 12'h777;
      20'h0b110: out <= 12'h000;
      20'h0b111: out <= 12'h000;
      20'h0b112: out <= 12'h000;
      20'h0b113: out <= 12'h000;
      20'h0b114: out <= 12'h000;
      20'h0b115: out <= 12'h000;
      20'h0b116: out <= 12'h000;
      20'h0b117: out <= 12'h000;
      20'h0b118: out <= 12'h000;
      20'h0b119: out <= 12'h000;
      20'h0b11a: out <= 12'h000;
      20'h0b11b: out <= 12'h000;
      20'h0b11c: out <= 12'h000;
      20'h0b11d: out <= 12'h000;
      20'h0b11e: out <= 12'h000;
      20'h0b11f: out <= 12'h000;
      20'h0b120: out <= 12'h000;
      20'h0b121: out <= 12'h000;
      20'h0b122: out <= 12'h000;
      20'h0b123: out <= 12'h000;
      20'h0b124: out <= 12'h000;
      20'h0b125: out <= 12'h000;
      20'h0b126: out <= 12'h000;
      20'h0b127: out <= 12'h000;
      20'h0b128: out <= 12'h000;
      20'h0b129: out <= 12'h000;
      20'h0b12a: out <= 12'h000;
      20'h0b12b: out <= 12'h000;
      20'h0b12c: out <= 12'h000;
      20'h0b12d: out <= 12'h000;
      20'h0b12e: out <= 12'h000;
      20'h0b12f: out <= 12'h000;
      20'h0b130: out <= 12'h088;
      20'h0b131: out <= 12'h088;
      20'h0b132: out <= 12'h088;
      20'h0b133: out <= 12'h088;
      20'h0b134: out <= 12'h088;
      20'h0b135: out <= 12'h088;
      20'h0b136: out <= 12'h088;
      20'h0b137: out <= 12'h088;
      20'h0b138: out <= 12'h088;
      20'h0b139: out <= 12'h088;
      20'h0b13a: out <= 12'h088;
      20'h0b13b: out <= 12'h088;
      20'h0b13c: out <= 12'h088;
      20'h0b13d: out <= 12'h088;
      20'h0b13e: out <= 12'h088;
      20'h0b13f: out <= 12'h088;
      20'h0b140: out <= 12'h088;
      20'h0b141: out <= 12'h088;
      20'h0b142: out <= 12'h088;
      20'h0b143: out <= 12'h088;
      20'h0b144: out <= 12'h088;
      20'h0b145: out <= 12'h088;
      20'h0b146: out <= 12'h088;
      20'h0b147: out <= 12'h088;
      20'h0b148: out <= 12'h088;
      20'h0b149: out <= 12'h088;
      20'h0b14a: out <= 12'h088;
      20'h0b14b: out <= 12'h088;
      20'h0b14c: out <= 12'h088;
      20'h0b14d: out <= 12'h088;
      20'h0b14e: out <= 12'h088;
      20'h0b14f: out <= 12'h088;
      20'h0b150: out <= 12'h088;
      20'h0b151: out <= 12'h088;
      20'h0b152: out <= 12'h088;
      20'h0b153: out <= 12'h088;
      20'h0b154: out <= 12'h088;
      20'h0b155: out <= 12'h088;
      20'h0b156: out <= 12'h088;
      20'h0b157: out <= 12'h088;
      20'h0b158: out <= 12'h088;
      20'h0b159: out <= 12'h088;
      20'h0b15a: out <= 12'h088;
      20'h0b15b: out <= 12'h088;
      20'h0b15c: out <= 12'h088;
      20'h0b15d: out <= 12'h088;
      20'h0b15e: out <= 12'h088;
      20'h0b15f: out <= 12'h088;
      20'h0b160: out <= 12'h088;
      20'h0b161: out <= 12'h088;
      20'h0b162: out <= 12'h088;
      20'h0b163: out <= 12'h088;
      20'h0b164: out <= 12'h088;
      20'h0b165: out <= 12'h088;
      20'h0b166: out <= 12'h088;
      20'h0b167: out <= 12'h088;
      20'h0b168: out <= 12'h088;
      20'h0b169: out <= 12'h088;
      20'h0b16a: out <= 12'h088;
      20'h0b16b: out <= 12'h088;
      20'h0b16c: out <= 12'h088;
      20'h0b16d: out <= 12'h088;
      20'h0b16e: out <= 12'h088;
      20'h0b16f: out <= 12'h088;
      20'h0b170: out <= 12'h088;
      20'h0b171: out <= 12'h088;
      20'h0b172: out <= 12'h088;
      20'h0b173: out <= 12'h088;
      20'h0b174: out <= 12'h088;
      20'h0b175: out <= 12'h088;
      20'h0b176: out <= 12'h088;
      20'h0b177: out <= 12'h088;
      20'h0b178: out <= 12'h088;
      20'h0b179: out <= 12'h088;
      20'h0b17a: out <= 12'h088;
      20'h0b17b: out <= 12'h088;
      20'h0b17c: out <= 12'h088;
      20'h0b17d: out <= 12'h088;
      20'h0b17e: out <= 12'h088;
      20'h0b17f: out <= 12'h088;
      20'h0b180: out <= 12'h088;
      20'h0b181: out <= 12'h088;
      20'h0b182: out <= 12'h088;
      20'h0b183: out <= 12'h088;
      20'h0b184: out <= 12'h088;
      20'h0b185: out <= 12'h088;
      20'h0b186: out <= 12'h088;
      20'h0b187: out <= 12'h088;
      20'h0b188: out <= 12'h088;
      20'h0b189: out <= 12'h088;
      20'h0b18a: out <= 12'h088;
      20'h0b18b: out <= 12'h088;
      20'h0b18c: out <= 12'h088;
      20'h0b18d: out <= 12'h088;
      20'h0b18e: out <= 12'h088;
      20'h0b18f: out <= 12'h088;
      20'h0b190: out <= 12'h088;
      20'h0b191: out <= 12'h088;
      20'h0b192: out <= 12'h088;
      20'h0b193: out <= 12'h088;
      20'h0b194: out <= 12'h088;
      20'h0b195: out <= 12'h088;
      20'h0b196: out <= 12'h088;
      20'h0b197: out <= 12'h088;
      20'h0b198: out <= 12'h088;
      20'h0b199: out <= 12'h603;
      20'h0b19a: out <= 12'h603;
      20'h0b19b: out <= 12'h603;
      20'h0b19c: out <= 12'h603;
      20'h0b19d: out <= 12'h603;
      20'h0b19e: out <= 12'h603;
      20'h0b19f: out <= 12'h603;
      20'h0b1a0: out <= 12'h603;
      20'h0b1a1: out <= 12'h603;
      20'h0b1a2: out <= 12'h603;
      20'h0b1a3: out <= 12'h603;
      20'h0b1a4: out <= 12'h603;
      20'h0b1a5: out <= 12'h603;
      20'h0b1a6: out <= 12'h603;
      20'h0b1a7: out <= 12'h603;
      20'h0b1a8: out <= 12'h603;
      20'h0b1a9: out <= 12'h603;
      20'h0b1aa: out <= 12'h603;
      20'h0b1ab: out <= 12'h603;
      20'h0b1ac: out <= 12'h603;
      20'h0b1ad: out <= 12'h603;
      20'h0b1ae: out <= 12'h603;
      20'h0b1af: out <= 12'h603;
      20'h0b1b0: out <= 12'h603;
      20'h0b1b1: out <= 12'h603;
      20'h0b1b2: out <= 12'h603;
      20'h0b1b3: out <= 12'h603;
      20'h0b1b4: out <= 12'h8d0;
      20'h0b1b5: out <= 12'h8d0;
      20'h0b1b6: out <= 12'h000;
      20'h0b1b7: out <= 12'h000;
      20'h0b1b8: out <= 12'h8d0;
      20'h0b1b9: out <= 12'h8d0;
      20'h0b1ba: out <= 12'h8d0;
      20'h0b1bb: out <= 12'h000;
      20'h0b1bc: out <= 12'h000;
      20'h0b1bd: out <= 12'h000;
      20'h0b1be: out <= 12'h000;
      20'h0b1bf: out <= 12'h8d0;
      20'h0b1c0: out <= 12'h8d0;
      20'h0b1c1: out <= 12'h000;
      20'h0b1c2: out <= 12'h000;
      20'h0b1c3: out <= 12'h000;
      20'h0b1c4: out <= 12'h000;
      20'h0b1c5: out <= 12'h000;
      20'h0b1c6: out <= 12'h000;
      20'h0b1c7: out <= 12'h000;
      20'h0b1c8: out <= 12'h000;
      20'h0b1c9: out <= 12'h8d0;
      20'h0b1ca: out <= 12'h8d0;
      20'h0b1cb: out <= 12'h000;
      20'h0b1cc: out <= 12'h000;
      20'h0b1cd: out <= 12'h000;
      20'h0b1ce: out <= 12'h000;
      20'h0b1cf: out <= 12'h000;
      20'h0b1d0: out <= 12'h000;
      20'h0b1d1: out <= 12'h8d0;
      20'h0b1d2: out <= 12'h8d0;
      20'h0b1d3: out <= 12'h000;
      20'h0b1d4: out <= 12'h000;
      20'h0b1d5: out <= 12'h8d0;
      20'h0b1d6: out <= 12'h8d0;
      20'h0b1d7: out <= 12'h000;
      20'h0b1d8: out <= 12'h8d0;
      20'h0b1d9: out <= 12'h8d0;
      20'h0b1da: out <= 12'h000;
      20'h0b1db: out <= 12'h000;
      20'h0b1dc: out <= 12'h8d0;
      20'h0b1dd: out <= 12'h8d0;
      20'h0b1de: out <= 12'h8d0;
      20'h0b1df: out <= 12'h8d0;
      20'h0b1e0: out <= 12'h8d0;
      20'h0b1e1: out <= 12'h8d0;
      20'h0b1e2: out <= 12'h000;
      20'h0b1e3: out <= 12'h000;
      20'h0b1e4: out <= 12'h8d0;
      20'h0b1e5: out <= 12'h8d0;
      20'h0b1e6: out <= 12'h000;
      20'h0b1e7: out <= 12'h000;
      20'h0b1e8: out <= 12'h000;
      20'h0b1e9: out <= 12'h000;
      20'h0b1ea: out <= 12'h000;
      20'h0b1eb: out <= 12'h000;
      20'h0b1ec: out <= 12'h000;
      20'h0b1ed: out <= 12'h000;
      20'h0b1ee: out <= 12'h000;
      20'h0b1ef: out <= 12'h000;
      20'h0b1f0: out <= 12'h8d0;
      20'h0b1f1: out <= 12'h8d0;
      20'h0b1f2: out <= 12'h000;
      20'h0b1f3: out <= 12'h000;
      20'h0b1f4: out <= 12'h8d0;
      20'h0b1f5: out <= 12'h8d0;
      20'h0b1f6: out <= 12'h000;
      20'h0b1f7: out <= 12'h000;
      20'h0b1f8: out <= 12'h000;
      20'h0b1f9: out <= 12'h8d0;
      20'h0b1fa: out <= 12'h8d0;
      20'h0b1fb: out <= 12'h000;
      20'h0b1fc: out <= 12'h8d0;
      20'h0b1fd: out <= 12'h8d0;
      20'h0b1fe: out <= 12'h000;
      20'h0b1ff: out <= 12'h000;
      20'h0b200: out <= 12'h000;
      20'h0b201: out <= 12'h8d0;
      20'h0b202: out <= 12'h8d0;
      20'h0b203: out <= 12'h000;
      20'h0b204: out <= 12'h603;
      20'h0b205: out <= 12'h603;
      20'h0b206: out <= 12'h603;
      20'h0b207: out <= 12'h603;
      20'h0b208: out <= 12'hee9;
      20'h0b209: out <= 12'hf87;
      20'h0b20a: out <= 12'hee9;
      20'h0b20b: out <= 12'hee9;
      20'h0b20c: out <= 12'hee9;
      20'h0b20d: out <= 12'hb27;
      20'h0b20e: out <= 12'hf87;
      20'h0b20f: out <= 12'hb27;
      20'h0b210: out <= 12'h000;
      20'h0b211: out <= 12'h000;
      20'h0b212: out <= 12'h000;
      20'h0b213: out <= 12'h000;
      20'h0b214: out <= 12'h000;
      20'h0b215: out <= 12'h000;
      20'h0b216: out <= 12'h000;
      20'h0b217: out <= 12'h000;
      20'h0b218: out <= 12'h777;
      20'h0b219: out <= 12'h555;
      20'h0b21a: out <= 12'h555;
      20'h0b21b: out <= 12'h555;
      20'h0b21c: out <= 12'h555;
      20'h0b21d: out <= 12'h555;
      20'h0b21e: out <= 12'h555;
      20'h0b21f: out <= 12'h555;
      20'h0b220: out <= 12'h555;
      20'h0b221: out <= 12'h555;
      20'h0b222: out <= 12'h555;
      20'h0b223: out <= 12'h555;
      20'h0b224: out <= 12'h555;
      20'h0b225: out <= 12'h555;
      20'h0b226: out <= 12'h555;
      20'h0b227: out <= 12'h777;
      20'h0b228: out <= 12'h000;
      20'h0b229: out <= 12'h000;
      20'h0b22a: out <= 12'h000;
      20'h0b22b: out <= 12'h000;
      20'h0b22c: out <= 12'h000;
      20'h0b22d: out <= 12'h000;
      20'h0b22e: out <= 12'h000;
      20'h0b22f: out <= 12'h000;
      20'h0b230: out <= 12'h000;
      20'h0b231: out <= 12'h000;
      20'h0b232: out <= 12'h000;
      20'h0b233: out <= 12'h000;
      20'h0b234: out <= 12'h000;
      20'h0b235: out <= 12'h000;
      20'h0b236: out <= 12'h000;
      20'h0b237: out <= 12'h000;
      20'h0b238: out <= 12'h000;
      20'h0b239: out <= 12'h000;
      20'h0b23a: out <= 12'h000;
      20'h0b23b: out <= 12'h000;
      20'h0b23c: out <= 12'h000;
      20'h0b23d: out <= 12'h000;
      20'h0b23e: out <= 12'h000;
      20'h0b23f: out <= 12'h000;
      20'h0b240: out <= 12'h000;
      20'h0b241: out <= 12'h000;
      20'h0b242: out <= 12'h000;
      20'h0b243: out <= 12'h000;
      20'h0b244: out <= 12'h000;
      20'h0b245: out <= 12'h000;
      20'h0b246: out <= 12'h000;
      20'h0b247: out <= 12'h000;
      20'h0b248: out <= 12'h088;
      20'h0b249: out <= 12'h088;
      20'h0b24a: out <= 12'h088;
      20'h0b24b: out <= 12'h088;
      20'h0b24c: out <= 12'h088;
      20'h0b24d: out <= 12'h088;
      20'h0b24e: out <= 12'h088;
      20'h0b24f: out <= 12'h088;
      20'h0b250: out <= 12'h088;
      20'h0b251: out <= 12'h088;
      20'h0b252: out <= 12'h088;
      20'h0b253: out <= 12'h088;
      20'h0b254: out <= 12'h088;
      20'h0b255: out <= 12'h088;
      20'h0b256: out <= 12'h088;
      20'h0b257: out <= 12'h088;
      20'h0b258: out <= 12'h088;
      20'h0b259: out <= 12'h088;
      20'h0b25a: out <= 12'h088;
      20'h0b25b: out <= 12'h088;
      20'h0b25c: out <= 12'h088;
      20'h0b25d: out <= 12'h088;
      20'h0b25e: out <= 12'h088;
      20'h0b25f: out <= 12'h088;
      20'h0b260: out <= 12'h088;
      20'h0b261: out <= 12'h088;
      20'h0b262: out <= 12'h088;
      20'h0b263: out <= 12'h088;
      20'h0b264: out <= 12'h088;
      20'h0b265: out <= 12'h088;
      20'h0b266: out <= 12'h088;
      20'h0b267: out <= 12'h088;
      20'h0b268: out <= 12'h088;
      20'h0b269: out <= 12'h088;
      20'h0b26a: out <= 12'h088;
      20'h0b26b: out <= 12'h088;
      20'h0b26c: out <= 12'h088;
      20'h0b26d: out <= 12'h088;
      20'h0b26e: out <= 12'h088;
      20'h0b26f: out <= 12'h088;
      20'h0b270: out <= 12'h088;
      20'h0b271: out <= 12'h088;
      20'h0b272: out <= 12'h088;
      20'h0b273: out <= 12'h088;
      20'h0b274: out <= 12'h088;
      20'h0b275: out <= 12'h088;
      20'h0b276: out <= 12'h088;
      20'h0b277: out <= 12'h088;
      20'h0b278: out <= 12'h088;
      20'h0b279: out <= 12'h088;
      20'h0b27a: out <= 12'h088;
      20'h0b27b: out <= 12'h088;
      20'h0b27c: out <= 12'h088;
      20'h0b27d: out <= 12'h088;
      20'h0b27e: out <= 12'h088;
      20'h0b27f: out <= 12'h088;
      20'h0b280: out <= 12'h088;
      20'h0b281: out <= 12'h088;
      20'h0b282: out <= 12'h088;
      20'h0b283: out <= 12'h088;
      20'h0b284: out <= 12'h088;
      20'h0b285: out <= 12'h088;
      20'h0b286: out <= 12'h088;
      20'h0b287: out <= 12'h088;
      20'h0b288: out <= 12'h088;
      20'h0b289: out <= 12'h088;
      20'h0b28a: out <= 12'h088;
      20'h0b28b: out <= 12'h088;
      20'h0b28c: out <= 12'h088;
      20'h0b28d: out <= 12'h088;
      20'h0b28e: out <= 12'h088;
      20'h0b28f: out <= 12'h088;
      20'h0b290: out <= 12'h088;
      20'h0b291: out <= 12'h088;
      20'h0b292: out <= 12'h088;
      20'h0b293: out <= 12'h088;
      20'h0b294: out <= 12'h088;
      20'h0b295: out <= 12'h088;
      20'h0b296: out <= 12'h088;
      20'h0b297: out <= 12'h088;
      20'h0b298: out <= 12'h088;
      20'h0b299: out <= 12'h088;
      20'h0b29a: out <= 12'h088;
      20'h0b29b: out <= 12'h088;
      20'h0b29c: out <= 12'h088;
      20'h0b29d: out <= 12'h088;
      20'h0b29e: out <= 12'h088;
      20'h0b29f: out <= 12'h088;
      20'h0b2a0: out <= 12'h088;
      20'h0b2a1: out <= 12'h088;
      20'h0b2a2: out <= 12'h088;
      20'h0b2a3: out <= 12'h088;
      20'h0b2a4: out <= 12'h088;
      20'h0b2a5: out <= 12'h088;
      20'h0b2a6: out <= 12'h088;
      20'h0b2a7: out <= 12'h088;
      20'h0b2a8: out <= 12'h088;
      20'h0b2a9: out <= 12'h088;
      20'h0b2aa: out <= 12'h088;
      20'h0b2ab: out <= 12'h088;
      20'h0b2ac: out <= 12'h088;
      20'h0b2ad: out <= 12'h088;
      20'h0b2ae: out <= 12'h088;
      20'h0b2af: out <= 12'h088;
      20'h0b2b0: out <= 12'h088;
      20'h0b2b1: out <= 12'h603;
      20'h0b2b2: out <= 12'h603;
      20'h0b2b3: out <= 12'h603;
      20'h0b2b4: out <= 12'h603;
      20'h0b2b5: out <= 12'h603;
      20'h0b2b6: out <= 12'h603;
      20'h0b2b7: out <= 12'h603;
      20'h0b2b8: out <= 12'h603;
      20'h0b2b9: out <= 12'h603;
      20'h0b2ba: out <= 12'h603;
      20'h0b2bb: out <= 12'h603;
      20'h0b2bc: out <= 12'h603;
      20'h0b2bd: out <= 12'h603;
      20'h0b2be: out <= 12'h603;
      20'h0b2bf: out <= 12'h603;
      20'h0b2c0: out <= 12'h603;
      20'h0b2c1: out <= 12'h603;
      20'h0b2c2: out <= 12'h603;
      20'h0b2c3: out <= 12'h603;
      20'h0b2c4: out <= 12'h603;
      20'h0b2c5: out <= 12'h603;
      20'h0b2c6: out <= 12'h603;
      20'h0b2c7: out <= 12'h603;
      20'h0b2c8: out <= 12'h603;
      20'h0b2c9: out <= 12'h603;
      20'h0b2ca: out <= 12'h603;
      20'h0b2cb: out <= 12'h603;
      20'h0b2cc: out <= 12'h8d0;
      20'h0b2cd: out <= 12'h8d0;
      20'h0b2ce: out <= 12'h000;
      20'h0b2cf: out <= 12'h8d0;
      20'h0b2d0: out <= 12'h000;
      20'h0b2d1: out <= 12'h8d0;
      20'h0b2d2: out <= 12'h8d0;
      20'h0b2d3: out <= 12'h000;
      20'h0b2d4: out <= 12'h000;
      20'h0b2d5: out <= 12'h000;
      20'h0b2d6: out <= 12'h000;
      20'h0b2d7: out <= 12'h8d0;
      20'h0b2d8: out <= 12'h8d0;
      20'h0b2d9: out <= 12'h000;
      20'h0b2da: out <= 12'h000;
      20'h0b2db: out <= 12'h000;
      20'h0b2dc: out <= 12'h000;
      20'h0b2dd: out <= 12'h000;
      20'h0b2de: out <= 12'h000;
      20'h0b2df: out <= 12'h8d0;
      20'h0b2e0: out <= 12'h8d0;
      20'h0b2e1: out <= 12'h8d0;
      20'h0b2e2: out <= 12'h000;
      20'h0b2e3: out <= 12'h000;
      20'h0b2e4: out <= 12'h000;
      20'h0b2e5: out <= 12'h000;
      20'h0b2e6: out <= 12'h8d0;
      20'h0b2e7: out <= 12'h8d0;
      20'h0b2e8: out <= 12'h8d0;
      20'h0b2e9: out <= 12'h8d0;
      20'h0b2ea: out <= 12'h000;
      20'h0b2eb: out <= 12'h000;
      20'h0b2ec: out <= 12'h8d0;
      20'h0b2ed: out <= 12'h8d0;
      20'h0b2ee: out <= 12'h000;
      20'h0b2ef: out <= 12'h000;
      20'h0b2f0: out <= 12'h8d0;
      20'h0b2f1: out <= 12'h8d0;
      20'h0b2f2: out <= 12'h000;
      20'h0b2f3: out <= 12'h000;
      20'h0b2f4: out <= 12'h000;
      20'h0b2f5: out <= 12'h000;
      20'h0b2f6: out <= 12'h000;
      20'h0b2f7: out <= 12'h000;
      20'h0b2f8: out <= 12'h000;
      20'h0b2f9: out <= 12'h8d0;
      20'h0b2fa: out <= 12'h8d0;
      20'h0b2fb: out <= 12'h000;
      20'h0b2fc: out <= 12'h8d0;
      20'h0b2fd: out <= 12'h8d0;
      20'h0b2fe: out <= 12'h8d0;
      20'h0b2ff: out <= 12'h8d0;
      20'h0b300: out <= 12'h8d0;
      20'h0b301: out <= 12'h8d0;
      20'h0b302: out <= 12'h000;
      20'h0b303: out <= 12'h000;
      20'h0b304: out <= 12'h000;
      20'h0b305: out <= 12'h000;
      20'h0b306: out <= 12'h000;
      20'h0b307: out <= 12'h8d0;
      20'h0b308: out <= 12'h8d0;
      20'h0b309: out <= 12'h000;
      20'h0b30a: out <= 12'h000;
      20'h0b30b: out <= 12'h000;
      20'h0b30c: out <= 12'h000;
      20'h0b30d: out <= 12'h8d0;
      20'h0b30e: out <= 12'h8d0;
      20'h0b30f: out <= 12'h8d0;
      20'h0b310: out <= 12'h8d0;
      20'h0b311: out <= 12'h8d0;
      20'h0b312: out <= 12'h000;
      20'h0b313: out <= 12'h000;
      20'h0b314: out <= 12'h000;
      20'h0b315: out <= 12'h8d0;
      20'h0b316: out <= 12'h8d0;
      20'h0b317: out <= 12'h8d0;
      20'h0b318: out <= 12'h8d0;
      20'h0b319: out <= 12'h8d0;
      20'h0b31a: out <= 12'h8d0;
      20'h0b31b: out <= 12'h000;
      20'h0b31c: out <= 12'h603;
      20'h0b31d: out <= 12'h603;
      20'h0b31e: out <= 12'h603;
      20'h0b31f: out <= 12'h603;
      20'h0b320: out <= 12'hee9;
      20'h0b321: out <= 12'hf87;
      20'h0b322: out <= 12'hee9;
      20'h0b323: out <= 12'hf87;
      20'h0b324: out <= 12'hf87;
      20'h0b325: out <= 12'hb27;
      20'h0b326: out <= 12'hf87;
      20'h0b327: out <= 12'hb27;
      20'h0b328: out <= 12'h000;
      20'h0b329: out <= 12'h000;
      20'h0b32a: out <= 12'h000;
      20'h0b32b: out <= 12'h000;
      20'h0b32c: out <= 12'h000;
      20'h0b32d: out <= 12'h000;
      20'h0b32e: out <= 12'h000;
      20'h0b32f: out <= 12'h000;
      20'h0b330: out <= 12'h777;
      20'h0b331: out <= 12'h555;
      20'h0b332: out <= 12'h555;
      20'h0b333: out <= 12'h555;
      20'h0b334: out <= 12'h555;
      20'h0b335: out <= 12'h555;
      20'h0b336: out <= 12'h555;
      20'h0b337: out <= 12'h555;
      20'h0b338: out <= 12'h555;
      20'h0b339: out <= 12'h555;
      20'h0b33a: out <= 12'h555;
      20'h0b33b: out <= 12'h555;
      20'h0b33c: out <= 12'h555;
      20'h0b33d: out <= 12'h555;
      20'h0b33e: out <= 12'h555;
      20'h0b33f: out <= 12'h777;
      20'h0b340: out <= 12'h000;
      20'h0b341: out <= 12'h000;
      20'h0b342: out <= 12'h000;
      20'h0b343: out <= 12'h000;
      20'h0b344: out <= 12'h000;
      20'h0b345: out <= 12'h000;
      20'h0b346: out <= 12'h000;
      20'h0b347: out <= 12'h000;
      20'h0b348: out <= 12'h000;
      20'h0b349: out <= 12'h000;
      20'h0b34a: out <= 12'h000;
      20'h0b34b: out <= 12'h000;
      20'h0b34c: out <= 12'h000;
      20'h0b34d: out <= 12'h000;
      20'h0b34e: out <= 12'h000;
      20'h0b34f: out <= 12'h000;
      20'h0b350: out <= 12'h000;
      20'h0b351: out <= 12'h000;
      20'h0b352: out <= 12'h000;
      20'h0b353: out <= 12'h000;
      20'h0b354: out <= 12'h000;
      20'h0b355: out <= 12'h000;
      20'h0b356: out <= 12'h000;
      20'h0b357: out <= 12'h000;
      20'h0b358: out <= 12'h000;
      20'h0b359: out <= 12'h000;
      20'h0b35a: out <= 12'h000;
      20'h0b35b: out <= 12'h000;
      20'h0b35c: out <= 12'h000;
      20'h0b35d: out <= 12'h000;
      20'h0b35e: out <= 12'h000;
      20'h0b35f: out <= 12'h000;
      20'h0b360: out <= 12'h088;
      20'h0b361: out <= 12'h088;
      20'h0b362: out <= 12'h088;
      20'h0b363: out <= 12'h088;
      20'h0b364: out <= 12'h088;
      20'h0b365: out <= 12'h088;
      20'h0b366: out <= 12'h088;
      20'h0b367: out <= 12'h088;
      20'h0b368: out <= 12'h088;
      20'h0b369: out <= 12'h088;
      20'h0b36a: out <= 12'h088;
      20'h0b36b: out <= 12'h088;
      20'h0b36c: out <= 12'h088;
      20'h0b36d: out <= 12'h088;
      20'h0b36e: out <= 12'h088;
      20'h0b36f: out <= 12'h088;
      20'h0b370: out <= 12'h088;
      20'h0b371: out <= 12'h088;
      20'h0b372: out <= 12'h088;
      20'h0b373: out <= 12'h088;
      20'h0b374: out <= 12'h088;
      20'h0b375: out <= 12'h088;
      20'h0b376: out <= 12'h088;
      20'h0b377: out <= 12'h088;
      20'h0b378: out <= 12'h088;
      20'h0b379: out <= 12'h088;
      20'h0b37a: out <= 12'h088;
      20'h0b37b: out <= 12'h088;
      20'h0b37c: out <= 12'h088;
      20'h0b37d: out <= 12'h088;
      20'h0b37e: out <= 12'h088;
      20'h0b37f: out <= 12'h088;
      20'h0b380: out <= 12'h088;
      20'h0b381: out <= 12'h088;
      20'h0b382: out <= 12'h088;
      20'h0b383: out <= 12'h088;
      20'h0b384: out <= 12'h088;
      20'h0b385: out <= 12'h088;
      20'h0b386: out <= 12'h088;
      20'h0b387: out <= 12'h088;
      20'h0b388: out <= 12'h088;
      20'h0b389: out <= 12'h088;
      20'h0b38a: out <= 12'h088;
      20'h0b38b: out <= 12'h088;
      20'h0b38c: out <= 12'h088;
      20'h0b38d: out <= 12'h088;
      20'h0b38e: out <= 12'h088;
      20'h0b38f: out <= 12'h088;
      20'h0b390: out <= 12'h088;
      20'h0b391: out <= 12'h088;
      20'h0b392: out <= 12'h088;
      20'h0b393: out <= 12'h088;
      20'h0b394: out <= 12'h088;
      20'h0b395: out <= 12'h088;
      20'h0b396: out <= 12'h088;
      20'h0b397: out <= 12'h088;
      20'h0b398: out <= 12'h088;
      20'h0b399: out <= 12'h088;
      20'h0b39a: out <= 12'h088;
      20'h0b39b: out <= 12'h088;
      20'h0b39c: out <= 12'h088;
      20'h0b39d: out <= 12'h088;
      20'h0b39e: out <= 12'h088;
      20'h0b39f: out <= 12'h088;
      20'h0b3a0: out <= 12'h088;
      20'h0b3a1: out <= 12'h088;
      20'h0b3a2: out <= 12'h088;
      20'h0b3a3: out <= 12'h088;
      20'h0b3a4: out <= 12'h088;
      20'h0b3a5: out <= 12'h088;
      20'h0b3a6: out <= 12'h088;
      20'h0b3a7: out <= 12'h088;
      20'h0b3a8: out <= 12'h088;
      20'h0b3a9: out <= 12'h088;
      20'h0b3aa: out <= 12'h088;
      20'h0b3ab: out <= 12'h088;
      20'h0b3ac: out <= 12'h088;
      20'h0b3ad: out <= 12'h088;
      20'h0b3ae: out <= 12'h088;
      20'h0b3af: out <= 12'h088;
      20'h0b3b0: out <= 12'h088;
      20'h0b3b1: out <= 12'h088;
      20'h0b3b2: out <= 12'h088;
      20'h0b3b3: out <= 12'h088;
      20'h0b3b4: out <= 12'h088;
      20'h0b3b5: out <= 12'h088;
      20'h0b3b6: out <= 12'h088;
      20'h0b3b7: out <= 12'h088;
      20'h0b3b8: out <= 12'h088;
      20'h0b3b9: out <= 12'h088;
      20'h0b3ba: out <= 12'h088;
      20'h0b3bb: out <= 12'h088;
      20'h0b3bc: out <= 12'h088;
      20'h0b3bd: out <= 12'h088;
      20'h0b3be: out <= 12'h088;
      20'h0b3bf: out <= 12'h088;
      20'h0b3c0: out <= 12'h088;
      20'h0b3c1: out <= 12'h088;
      20'h0b3c2: out <= 12'h088;
      20'h0b3c3: out <= 12'h088;
      20'h0b3c4: out <= 12'h088;
      20'h0b3c5: out <= 12'h088;
      20'h0b3c6: out <= 12'h088;
      20'h0b3c7: out <= 12'h088;
      20'h0b3c8: out <= 12'h088;
      20'h0b3c9: out <= 12'h222;
      20'h0b3ca: out <= 12'h222;
      20'h0b3cb: out <= 12'h222;
      20'h0b3cc: out <= 12'h222;
      20'h0b3cd: out <= 12'h222;
      20'h0b3ce: out <= 12'h222;
      20'h0b3cf: out <= 12'h222;
      20'h0b3d0: out <= 12'h222;
      20'h0b3d1: out <= 12'h222;
      20'h0b3d2: out <= 12'h222;
      20'h0b3d3: out <= 12'h222;
      20'h0b3d4: out <= 12'h222;
      20'h0b3d5: out <= 12'h222;
      20'h0b3d6: out <= 12'h222;
      20'h0b3d7: out <= 12'h222;
      20'h0b3d8: out <= 12'h222;
      20'h0b3d9: out <= 12'h222;
      20'h0b3da: out <= 12'h222;
      20'h0b3db: out <= 12'h222;
      20'h0b3dc: out <= 12'h222;
      20'h0b3dd: out <= 12'h222;
      20'h0b3de: out <= 12'h222;
      20'h0b3df: out <= 12'h222;
      20'h0b3e0: out <= 12'h603;
      20'h0b3e1: out <= 12'h603;
      20'h0b3e2: out <= 12'h603;
      20'h0b3e3: out <= 12'h603;
      20'h0b3e4: out <= 12'h8d0;
      20'h0b3e5: out <= 12'h8d0;
      20'h0b3e6: out <= 12'h8d0;
      20'h0b3e7: out <= 12'h000;
      20'h0b3e8: out <= 12'h000;
      20'h0b3e9: out <= 12'h8d0;
      20'h0b3ea: out <= 12'h8d0;
      20'h0b3eb: out <= 12'h000;
      20'h0b3ec: out <= 12'h000;
      20'h0b3ed: out <= 12'h000;
      20'h0b3ee: out <= 12'h000;
      20'h0b3ef: out <= 12'h8d0;
      20'h0b3f0: out <= 12'h8d0;
      20'h0b3f1: out <= 12'h000;
      20'h0b3f2: out <= 12'h000;
      20'h0b3f3: out <= 12'h000;
      20'h0b3f4: out <= 12'h000;
      20'h0b3f5: out <= 12'h8d0;
      20'h0b3f6: out <= 12'h8d0;
      20'h0b3f7: out <= 12'h8d0;
      20'h0b3f8: out <= 12'h000;
      20'h0b3f9: out <= 12'h000;
      20'h0b3fa: out <= 12'h000;
      20'h0b3fb: out <= 12'h000;
      20'h0b3fc: out <= 12'h000;
      20'h0b3fd: out <= 12'h000;
      20'h0b3fe: out <= 12'h000;
      20'h0b3ff: out <= 12'h000;
      20'h0b400: out <= 12'h000;
      20'h0b401: out <= 12'h8d0;
      20'h0b402: out <= 12'h8d0;
      20'h0b403: out <= 12'h000;
      20'h0b404: out <= 12'h8d0;
      20'h0b405: out <= 12'h8d0;
      20'h0b406: out <= 12'h8d0;
      20'h0b407: out <= 12'h8d0;
      20'h0b408: out <= 12'h8d0;
      20'h0b409: out <= 12'h8d0;
      20'h0b40a: out <= 12'h8d0;
      20'h0b40b: out <= 12'h000;
      20'h0b40c: out <= 12'h000;
      20'h0b40d: out <= 12'h000;
      20'h0b40e: out <= 12'h000;
      20'h0b40f: out <= 12'h000;
      20'h0b410: out <= 12'h000;
      20'h0b411: out <= 12'h8d0;
      20'h0b412: out <= 12'h8d0;
      20'h0b413: out <= 12'h000;
      20'h0b414: out <= 12'h8d0;
      20'h0b415: out <= 12'h8d0;
      20'h0b416: out <= 12'h000;
      20'h0b417: out <= 12'h000;
      20'h0b418: out <= 12'h000;
      20'h0b419: out <= 12'h8d0;
      20'h0b41a: out <= 12'h8d0;
      20'h0b41b: out <= 12'h000;
      20'h0b41c: out <= 12'h000;
      20'h0b41d: out <= 12'h000;
      20'h0b41e: out <= 12'h8d0;
      20'h0b41f: out <= 12'h8d0;
      20'h0b420: out <= 12'h000;
      20'h0b421: out <= 12'h000;
      20'h0b422: out <= 12'h000;
      20'h0b423: out <= 12'h000;
      20'h0b424: out <= 12'h8d0;
      20'h0b425: out <= 12'h8d0;
      20'h0b426: out <= 12'h000;
      20'h0b427: out <= 12'h000;
      20'h0b428: out <= 12'h000;
      20'h0b429: out <= 12'h8d0;
      20'h0b42a: out <= 12'h8d0;
      20'h0b42b: out <= 12'h000;
      20'h0b42c: out <= 12'h000;
      20'h0b42d: out <= 12'h000;
      20'h0b42e: out <= 12'h000;
      20'h0b42f: out <= 12'h000;
      20'h0b430: out <= 12'h000;
      20'h0b431: out <= 12'h8d0;
      20'h0b432: out <= 12'h8d0;
      20'h0b433: out <= 12'h000;
      20'h0b434: out <= 12'h603;
      20'h0b435: out <= 12'h603;
      20'h0b436: out <= 12'h603;
      20'h0b437: out <= 12'h603;
      20'h0b438: out <= 12'hee9;
      20'h0b439: out <= 12'hf87;
      20'h0b43a: out <= 12'hee9;
      20'h0b43b: out <= 12'hf87;
      20'h0b43c: out <= 12'hf87;
      20'h0b43d: out <= 12'hb27;
      20'h0b43e: out <= 12'hf87;
      20'h0b43f: out <= 12'hb27;
      20'h0b440: out <= 12'h000;
      20'h0b441: out <= 12'h000;
      20'h0b442: out <= 12'h000;
      20'h0b443: out <= 12'h000;
      20'h0b444: out <= 12'h000;
      20'h0b445: out <= 12'h000;
      20'h0b446: out <= 12'h000;
      20'h0b447: out <= 12'h000;
      20'h0b448: out <= 12'h777;
      20'h0b449: out <= 12'h555;
      20'h0b44a: out <= 12'h555;
      20'h0b44b: out <= 12'h555;
      20'h0b44c: out <= 12'h555;
      20'h0b44d: out <= 12'h555;
      20'h0b44e: out <= 12'h555;
      20'h0b44f: out <= 12'h555;
      20'h0b450: out <= 12'h555;
      20'h0b451: out <= 12'h555;
      20'h0b452: out <= 12'h555;
      20'h0b453: out <= 12'h555;
      20'h0b454: out <= 12'h555;
      20'h0b455: out <= 12'h555;
      20'h0b456: out <= 12'h555;
      20'h0b457: out <= 12'h777;
      20'h0b458: out <= 12'h000;
      20'h0b459: out <= 12'h000;
      20'h0b45a: out <= 12'h000;
      20'h0b45b: out <= 12'h000;
      20'h0b45c: out <= 12'h000;
      20'h0b45d: out <= 12'h000;
      20'h0b45e: out <= 12'h000;
      20'h0b45f: out <= 12'h000;
      20'h0b460: out <= 12'h000;
      20'h0b461: out <= 12'h000;
      20'h0b462: out <= 12'h000;
      20'h0b463: out <= 12'h000;
      20'h0b464: out <= 12'h000;
      20'h0b465: out <= 12'h000;
      20'h0b466: out <= 12'h000;
      20'h0b467: out <= 12'h000;
      20'h0b468: out <= 12'h000;
      20'h0b469: out <= 12'h000;
      20'h0b46a: out <= 12'h000;
      20'h0b46b: out <= 12'h000;
      20'h0b46c: out <= 12'h000;
      20'h0b46d: out <= 12'h000;
      20'h0b46e: out <= 12'h000;
      20'h0b46f: out <= 12'h000;
      20'h0b470: out <= 12'h000;
      20'h0b471: out <= 12'h000;
      20'h0b472: out <= 12'h000;
      20'h0b473: out <= 12'h000;
      20'h0b474: out <= 12'h000;
      20'h0b475: out <= 12'h000;
      20'h0b476: out <= 12'h000;
      20'h0b477: out <= 12'h000;
      20'h0b478: out <= 12'h088;
      20'h0b479: out <= 12'h088;
      20'h0b47a: out <= 12'h088;
      20'h0b47b: out <= 12'h088;
      20'h0b47c: out <= 12'h088;
      20'h0b47d: out <= 12'h088;
      20'h0b47e: out <= 12'h088;
      20'h0b47f: out <= 12'h088;
      20'h0b480: out <= 12'h088;
      20'h0b481: out <= 12'h088;
      20'h0b482: out <= 12'h088;
      20'h0b483: out <= 12'h088;
      20'h0b484: out <= 12'h088;
      20'h0b485: out <= 12'h088;
      20'h0b486: out <= 12'h088;
      20'h0b487: out <= 12'h088;
      20'h0b488: out <= 12'h088;
      20'h0b489: out <= 12'h088;
      20'h0b48a: out <= 12'h088;
      20'h0b48b: out <= 12'h088;
      20'h0b48c: out <= 12'h088;
      20'h0b48d: out <= 12'h088;
      20'h0b48e: out <= 12'h088;
      20'h0b48f: out <= 12'h088;
      20'h0b490: out <= 12'h088;
      20'h0b491: out <= 12'h088;
      20'h0b492: out <= 12'h088;
      20'h0b493: out <= 12'h088;
      20'h0b494: out <= 12'h088;
      20'h0b495: out <= 12'h088;
      20'h0b496: out <= 12'h088;
      20'h0b497: out <= 12'h088;
      20'h0b498: out <= 12'h088;
      20'h0b499: out <= 12'h088;
      20'h0b49a: out <= 12'h088;
      20'h0b49b: out <= 12'h088;
      20'h0b49c: out <= 12'h088;
      20'h0b49d: out <= 12'h088;
      20'h0b49e: out <= 12'h088;
      20'h0b49f: out <= 12'h088;
      20'h0b4a0: out <= 12'h088;
      20'h0b4a1: out <= 12'h088;
      20'h0b4a2: out <= 12'h088;
      20'h0b4a3: out <= 12'h088;
      20'h0b4a4: out <= 12'h088;
      20'h0b4a5: out <= 12'h088;
      20'h0b4a6: out <= 12'h088;
      20'h0b4a7: out <= 12'h088;
      20'h0b4a8: out <= 12'h088;
      20'h0b4a9: out <= 12'h088;
      20'h0b4aa: out <= 12'h088;
      20'h0b4ab: out <= 12'h088;
      20'h0b4ac: out <= 12'h088;
      20'h0b4ad: out <= 12'h088;
      20'h0b4ae: out <= 12'h088;
      20'h0b4af: out <= 12'h088;
      20'h0b4b0: out <= 12'h088;
      20'h0b4b1: out <= 12'h088;
      20'h0b4b2: out <= 12'h088;
      20'h0b4b3: out <= 12'h088;
      20'h0b4b4: out <= 12'h088;
      20'h0b4b5: out <= 12'h088;
      20'h0b4b6: out <= 12'h088;
      20'h0b4b7: out <= 12'h088;
      20'h0b4b8: out <= 12'h088;
      20'h0b4b9: out <= 12'h088;
      20'h0b4ba: out <= 12'h088;
      20'h0b4bb: out <= 12'h088;
      20'h0b4bc: out <= 12'h088;
      20'h0b4bd: out <= 12'h088;
      20'h0b4be: out <= 12'h088;
      20'h0b4bf: out <= 12'h088;
      20'h0b4c0: out <= 12'h088;
      20'h0b4c1: out <= 12'h088;
      20'h0b4c2: out <= 12'h088;
      20'h0b4c3: out <= 12'h088;
      20'h0b4c4: out <= 12'h088;
      20'h0b4c5: out <= 12'h088;
      20'h0b4c6: out <= 12'h088;
      20'h0b4c7: out <= 12'h088;
      20'h0b4c8: out <= 12'h088;
      20'h0b4c9: out <= 12'h088;
      20'h0b4ca: out <= 12'h088;
      20'h0b4cb: out <= 12'h088;
      20'h0b4cc: out <= 12'h088;
      20'h0b4cd: out <= 12'h088;
      20'h0b4ce: out <= 12'h088;
      20'h0b4cf: out <= 12'h088;
      20'h0b4d0: out <= 12'h088;
      20'h0b4d1: out <= 12'h088;
      20'h0b4d2: out <= 12'h088;
      20'h0b4d3: out <= 12'h088;
      20'h0b4d4: out <= 12'h088;
      20'h0b4d5: out <= 12'h088;
      20'h0b4d6: out <= 12'h088;
      20'h0b4d7: out <= 12'h088;
      20'h0b4d8: out <= 12'h088;
      20'h0b4d9: out <= 12'h088;
      20'h0b4da: out <= 12'h088;
      20'h0b4db: out <= 12'h088;
      20'h0b4dc: out <= 12'h088;
      20'h0b4dd: out <= 12'h088;
      20'h0b4de: out <= 12'h088;
      20'h0b4df: out <= 12'h088;
      20'h0b4e0: out <= 12'h088;
      20'h0b4e1: out <= 12'h222;
      20'h0b4e2: out <= 12'h222;
      20'h0b4e3: out <= 12'h222;
      20'h0b4e4: out <= 12'h222;
      20'h0b4e5: out <= 12'h222;
      20'h0b4e6: out <= 12'h222;
      20'h0b4e7: out <= 12'h222;
      20'h0b4e8: out <= 12'h222;
      20'h0b4e9: out <= 12'h222;
      20'h0b4ea: out <= 12'h222;
      20'h0b4eb: out <= 12'h222;
      20'h0b4ec: out <= 12'h222;
      20'h0b4ed: out <= 12'h222;
      20'h0b4ee: out <= 12'h222;
      20'h0b4ef: out <= 12'h222;
      20'h0b4f0: out <= 12'h222;
      20'h0b4f1: out <= 12'h222;
      20'h0b4f2: out <= 12'h222;
      20'h0b4f3: out <= 12'h222;
      20'h0b4f4: out <= 12'h222;
      20'h0b4f5: out <= 12'h222;
      20'h0b4f6: out <= 12'h222;
      20'h0b4f7: out <= 12'h222;
      20'h0b4f8: out <= 12'h603;
      20'h0b4f9: out <= 12'h603;
      20'h0b4fa: out <= 12'h603;
      20'h0b4fb: out <= 12'h603;
      20'h0b4fc: out <= 12'h8d0;
      20'h0b4fd: out <= 12'h8d0;
      20'h0b4fe: out <= 12'h000;
      20'h0b4ff: out <= 12'h000;
      20'h0b500: out <= 12'h000;
      20'h0b501: out <= 12'h8d0;
      20'h0b502: out <= 12'h8d0;
      20'h0b503: out <= 12'h000;
      20'h0b504: out <= 12'h000;
      20'h0b505: out <= 12'h000;
      20'h0b506: out <= 12'h000;
      20'h0b507: out <= 12'h8d0;
      20'h0b508: out <= 12'h8d0;
      20'h0b509: out <= 12'h000;
      20'h0b50a: out <= 12'h000;
      20'h0b50b: out <= 12'h000;
      20'h0b50c: out <= 12'h8d0;
      20'h0b50d: out <= 12'h8d0;
      20'h0b50e: out <= 12'h000;
      20'h0b50f: out <= 12'h000;
      20'h0b510: out <= 12'h000;
      20'h0b511: out <= 12'h000;
      20'h0b512: out <= 12'h000;
      20'h0b513: out <= 12'h000;
      20'h0b514: out <= 12'h8d0;
      20'h0b515: out <= 12'h8d0;
      20'h0b516: out <= 12'h000;
      20'h0b517: out <= 12'h000;
      20'h0b518: out <= 12'h000;
      20'h0b519: out <= 12'h8d0;
      20'h0b51a: out <= 12'h8d0;
      20'h0b51b: out <= 12'h000;
      20'h0b51c: out <= 12'h000;
      20'h0b51d: out <= 12'h000;
      20'h0b51e: out <= 12'h000;
      20'h0b51f: out <= 12'h000;
      20'h0b520: out <= 12'h8d0;
      20'h0b521: out <= 12'h8d0;
      20'h0b522: out <= 12'h000;
      20'h0b523: out <= 12'h000;
      20'h0b524: out <= 12'h8d0;
      20'h0b525: out <= 12'h8d0;
      20'h0b526: out <= 12'h000;
      20'h0b527: out <= 12'h000;
      20'h0b528: out <= 12'h000;
      20'h0b529: out <= 12'h8d0;
      20'h0b52a: out <= 12'h8d0;
      20'h0b52b: out <= 12'h000;
      20'h0b52c: out <= 12'h8d0;
      20'h0b52d: out <= 12'h8d0;
      20'h0b52e: out <= 12'h000;
      20'h0b52f: out <= 12'h000;
      20'h0b530: out <= 12'h000;
      20'h0b531: out <= 12'h8d0;
      20'h0b532: out <= 12'h8d0;
      20'h0b533: out <= 12'h000;
      20'h0b534: out <= 12'h000;
      20'h0b535: out <= 12'h000;
      20'h0b536: out <= 12'h8d0;
      20'h0b537: out <= 12'h8d0;
      20'h0b538: out <= 12'h000;
      20'h0b539: out <= 12'h000;
      20'h0b53a: out <= 12'h000;
      20'h0b53b: out <= 12'h000;
      20'h0b53c: out <= 12'h8d0;
      20'h0b53d: out <= 12'h8d0;
      20'h0b53e: out <= 12'h000;
      20'h0b53f: out <= 12'h000;
      20'h0b540: out <= 12'h000;
      20'h0b541: out <= 12'h8d0;
      20'h0b542: out <= 12'h8d0;
      20'h0b543: out <= 12'h000;
      20'h0b544: out <= 12'h000;
      20'h0b545: out <= 12'h000;
      20'h0b546: out <= 12'h000;
      20'h0b547: out <= 12'h000;
      20'h0b548: out <= 12'h8d0;
      20'h0b549: out <= 12'h8d0;
      20'h0b54a: out <= 12'h000;
      20'h0b54b: out <= 12'h000;
      20'h0b54c: out <= 12'h603;
      20'h0b54d: out <= 12'h603;
      20'h0b54e: out <= 12'h603;
      20'h0b54f: out <= 12'h603;
      20'h0b550: out <= 12'hee9;
      20'h0b551: out <= 12'hf87;
      20'h0b552: out <= 12'hee9;
      20'h0b553: out <= 12'hb27;
      20'h0b554: out <= 12'hb27;
      20'h0b555: out <= 12'hb27;
      20'h0b556: out <= 12'hf87;
      20'h0b557: out <= 12'hb27;
      20'h0b558: out <= 12'h000;
      20'h0b559: out <= 12'h000;
      20'h0b55a: out <= 12'h000;
      20'h0b55b: out <= 12'h000;
      20'h0b55c: out <= 12'h000;
      20'h0b55d: out <= 12'h000;
      20'h0b55e: out <= 12'h000;
      20'h0b55f: out <= 12'h000;
      20'h0b560: out <= 12'h777;
      20'h0b561: out <= 12'h555;
      20'h0b562: out <= 12'h555;
      20'h0b563: out <= 12'h555;
      20'h0b564: out <= 12'h555;
      20'h0b565: out <= 12'h555;
      20'h0b566: out <= 12'h555;
      20'h0b567: out <= 12'h555;
      20'h0b568: out <= 12'h555;
      20'h0b569: out <= 12'h555;
      20'h0b56a: out <= 12'h555;
      20'h0b56b: out <= 12'h555;
      20'h0b56c: out <= 12'h555;
      20'h0b56d: out <= 12'h555;
      20'h0b56e: out <= 12'h555;
      20'h0b56f: out <= 12'h777;
      20'h0b570: out <= 12'h000;
      20'h0b571: out <= 12'h000;
      20'h0b572: out <= 12'h000;
      20'h0b573: out <= 12'h000;
      20'h0b574: out <= 12'h000;
      20'h0b575: out <= 12'h000;
      20'h0b576: out <= 12'h000;
      20'h0b577: out <= 12'h000;
      20'h0b578: out <= 12'h000;
      20'h0b579: out <= 12'h000;
      20'h0b57a: out <= 12'h000;
      20'h0b57b: out <= 12'h000;
      20'h0b57c: out <= 12'h000;
      20'h0b57d: out <= 12'h000;
      20'h0b57e: out <= 12'h000;
      20'h0b57f: out <= 12'h000;
      20'h0b580: out <= 12'h000;
      20'h0b581: out <= 12'h000;
      20'h0b582: out <= 12'h000;
      20'h0b583: out <= 12'h000;
      20'h0b584: out <= 12'h000;
      20'h0b585: out <= 12'h000;
      20'h0b586: out <= 12'h000;
      20'h0b587: out <= 12'h000;
      20'h0b588: out <= 12'h000;
      20'h0b589: out <= 12'h000;
      20'h0b58a: out <= 12'h000;
      20'h0b58b: out <= 12'h000;
      20'h0b58c: out <= 12'h000;
      20'h0b58d: out <= 12'h000;
      20'h0b58e: out <= 12'h000;
      20'h0b58f: out <= 12'h000;
      20'h0b590: out <= 12'h088;
      20'h0b591: out <= 12'h088;
      20'h0b592: out <= 12'h088;
      20'h0b593: out <= 12'h088;
      20'h0b594: out <= 12'h088;
      20'h0b595: out <= 12'h088;
      20'h0b596: out <= 12'h088;
      20'h0b597: out <= 12'h088;
      20'h0b598: out <= 12'h088;
      20'h0b599: out <= 12'h088;
      20'h0b59a: out <= 12'h088;
      20'h0b59b: out <= 12'h088;
      20'h0b59c: out <= 12'h088;
      20'h0b59d: out <= 12'h088;
      20'h0b59e: out <= 12'h088;
      20'h0b59f: out <= 12'h088;
      20'h0b5a0: out <= 12'h088;
      20'h0b5a1: out <= 12'h088;
      20'h0b5a2: out <= 12'h088;
      20'h0b5a3: out <= 12'h088;
      20'h0b5a4: out <= 12'h088;
      20'h0b5a5: out <= 12'h088;
      20'h0b5a6: out <= 12'h088;
      20'h0b5a7: out <= 12'h088;
      20'h0b5a8: out <= 12'h088;
      20'h0b5a9: out <= 12'h088;
      20'h0b5aa: out <= 12'h088;
      20'h0b5ab: out <= 12'h088;
      20'h0b5ac: out <= 12'h088;
      20'h0b5ad: out <= 12'h088;
      20'h0b5ae: out <= 12'h088;
      20'h0b5af: out <= 12'h088;
      20'h0b5b0: out <= 12'h088;
      20'h0b5b1: out <= 12'h088;
      20'h0b5b2: out <= 12'h088;
      20'h0b5b3: out <= 12'h088;
      20'h0b5b4: out <= 12'h088;
      20'h0b5b5: out <= 12'h088;
      20'h0b5b6: out <= 12'h088;
      20'h0b5b7: out <= 12'h088;
      20'h0b5b8: out <= 12'h088;
      20'h0b5b9: out <= 12'h088;
      20'h0b5ba: out <= 12'h088;
      20'h0b5bb: out <= 12'h088;
      20'h0b5bc: out <= 12'h088;
      20'h0b5bd: out <= 12'h088;
      20'h0b5be: out <= 12'h088;
      20'h0b5bf: out <= 12'h088;
      20'h0b5c0: out <= 12'h088;
      20'h0b5c1: out <= 12'h088;
      20'h0b5c2: out <= 12'h088;
      20'h0b5c3: out <= 12'h088;
      20'h0b5c4: out <= 12'h088;
      20'h0b5c5: out <= 12'h088;
      20'h0b5c6: out <= 12'h088;
      20'h0b5c7: out <= 12'h088;
      20'h0b5c8: out <= 12'h088;
      20'h0b5c9: out <= 12'h088;
      20'h0b5ca: out <= 12'h088;
      20'h0b5cb: out <= 12'h088;
      20'h0b5cc: out <= 12'h088;
      20'h0b5cd: out <= 12'h088;
      20'h0b5ce: out <= 12'h088;
      20'h0b5cf: out <= 12'h088;
      20'h0b5d0: out <= 12'h088;
      20'h0b5d1: out <= 12'h088;
      20'h0b5d2: out <= 12'h088;
      20'h0b5d3: out <= 12'h088;
      20'h0b5d4: out <= 12'h088;
      20'h0b5d5: out <= 12'h088;
      20'h0b5d6: out <= 12'h088;
      20'h0b5d7: out <= 12'h088;
      20'h0b5d8: out <= 12'h088;
      20'h0b5d9: out <= 12'h088;
      20'h0b5da: out <= 12'h088;
      20'h0b5db: out <= 12'h088;
      20'h0b5dc: out <= 12'h088;
      20'h0b5dd: out <= 12'h088;
      20'h0b5de: out <= 12'h088;
      20'h0b5df: out <= 12'h088;
      20'h0b5e0: out <= 12'h088;
      20'h0b5e1: out <= 12'h088;
      20'h0b5e2: out <= 12'h088;
      20'h0b5e3: out <= 12'h088;
      20'h0b5e4: out <= 12'h088;
      20'h0b5e5: out <= 12'h088;
      20'h0b5e6: out <= 12'h088;
      20'h0b5e7: out <= 12'h088;
      20'h0b5e8: out <= 12'h088;
      20'h0b5e9: out <= 12'h088;
      20'h0b5ea: out <= 12'h088;
      20'h0b5eb: out <= 12'h088;
      20'h0b5ec: out <= 12'h088;
      20'h0b5ed: out <= 12'h088;
      20'h0b5ee: out <= 12'h088;
      20'h0b5ef: out <= 12'h088;
      20'h0b5f0: out <= 12'h088;
      20'h0b5f1: out <= 12'h088;
      20'h0b5f2: out <= 12'h088;
      20'h0b5f3: out <= 12'h088;
      20'h0b5f4: out <= 12'h088;
      20'h0b5f5: out <= 12'h088;
      20'h0b5f6: out <= 12'h088;
      20'h0b5f7: out <= 12'h088;
      20'h0b5f8: out <= 12'h088;
      20'h0b5f9: out <= 12'h222;
      20'h0b5fa: out <= 12'h222;
      20'h0b5fb: out <= 12'h222;
      20'h0b5fc: out <= 12'h222;
      20'h0b5fd: out <= 12'h222;
      20'h0b5fe: out <= 12'h222;
      20'h0b5ff: out <= 12'h222;
      20'h0b600: out <= 12'h222;
      20'h0b601: out <= 12'h222;
      20'h0b602: out <= 12'h222;
      20'h0b603: out <= 12'h222;
      20'h0b604: out <= 12'h660;
      20'h0b605: out <= 12'h222;
      20'h0b606: out <= 12'h222;
      20'h0b607: out <= 12'h222;
      20'h0b608: out <= 12'h222;
      20'h0b609: out <= 12'h222;
      20'h0b60a: out <= 12'h222;
      20'h0b60b: out <= 12'h222;
      20'h0b60c: out <= 12'h222;
      20'h0b60d: out <= 12'h222;
      20'h0b60e: out <= 12'h222;
      20'h0b60f: out <= 12'h222;
      20'h0b610: out <= 12'h603;
      20'h0b611: out <= 12'h603;
      20'h0b612: out <= 12'h603;
      20'h0b613: out <= 12'h603;
      20'h0b614: out <= 12'h000;
      20'h0b615: out <= 12'h8d0;
      20'h0b616: out <= 12'h8d0;
      20'h0b617: out <= 12'h8d0;
      20'h0b618: out <= 12'h8d0;
      20'h0b619: out <= 12'h8d0;
      20'h0b61a: out <= 12'h000;
      20'h0b61b: out <= 12'h000;
      20'h0b61c: out <= 12'h000;
      20'h0b61d: out <= 12'h000;
      20'h0b61e: out <= 12'h000;
      20'h0b61f: out <= 12'h8d0;
      20'h0b620: out <= 12'h8d0;
      20'h0b621: out <= 12'h000;
      20'h0b622: out <= 12'h000;
      20'h0b623: out <= 12'h000;
      20'h0b624: out <= 12'h8d0;
      20'h0b625: out <= 12'h8d0;
      20'h0b626: out <= 12'h8d0;
      20'h0b627: out <= 12'h8d0;
      20'h0b628: out <= 12'h8d0;
      20'h0b629: out <= 12'h8d0;
      20'h0b62a: out <= 12'h8d0;
      20'h0b62b: out <= 12'h000;
      20'h0b62c: out <= 12'h000;
      20'h0b62d: out <= 12'h8d0;
      20'h0b62e: out <= 12'h8d0;
      20'h0b62f: out <= 12'h8d0;
      20'h0b630: out <= 12'h8d0;
      20'h0b631: out <= 12'h8d0;
      20'h0b632: out <= 12'h000;
      20'h0b633: out <= 12'h000;
      20'h0b634: out <= 12'h000;
      20'h0b635: out <= 12'h000;
      20'h0b636: out <= 12'h000;
      20'h0b637: out <= 12'h000;
      20'h0b638: out <= 12'h8d0;
      20'h0b639: out <= 12'h8d0;
      20'h0b63a: out <= 12'h000;
      20'h0b63b: out <= 12'h000;
      20'h0b63c: out <= 12'h000;
      20'h0b63d: out <= 12'h8d0;
      20'h0b63e: out <= 12'h8d0;
      20'h0b63f: out <= 12'h8d0;
      20'h0b640: out <= 12'h8d0;
      20'h0b641: out <= 12'h8d0;
      20'h0b642: out <= 12'h000;
      20'h0b643: out <= 12'h000;
      20'h0b644: out <= 12'h000;
      20'h0b645: out <= 12'h8d0;
      20'h0b646: out <= 12'h8d0;
      20'h0b647: out <= 12'h8d0;
      20'h0b648: out <= 12'h8d0;
      20'h0b649: out <= 12'h8d0;
      20'h0b64a: out <= 12'h000;
      20'h0b64b: out <= 12'h000;
      20'h0b64c: out <= 12'h000;
      20'h0b64d: out <= 12'h000;
      20'h0b64e: out <= 12'h8d0;
      20'h0b64f: out <= 12'h8d0;
      20'h0b650: out <= 12'h000;
      20'h0b651: out <= 12'h000;
      20'h0b652: out <= 12'h000;
      20'h0b653: out <= 12'h000;
      20'h0b654: out <= 12'h000;
      20'h0b655: out <= 12'h8d0;
      20'h0b656: out <= 12'h8d0;
      20'h0b657: out <= 12'h8d0;
      20'h0b658: out <= 12'h8d0;
      20'h0b659: out <= 12'h8d0;
      20'h0b65a: out <= 12'h000;
      20'h0b65b: out <= 12'h000;
      20'h0b65c: out <= 12'h000;
      20'h0b65d: out <= 12'h8d0;
      20'h0b65e: out <= 12'h8d0;
      20'h0b65f: out <= 12'h8d0;
      20'h0b660: out <= 12'h8d0;
      20'h0b661: out <= 12'h000;
      20'h0b662: out <= 12'h000;
      20'h0b663: out <= 12'h000;
      20'h0b664: out <= 12'h603;
      20'h0b665: out <= 12'h603;
      20'h0b666: out <= 12'h603;
      20'h0b667: out <= 12'h603;
      20'h0b668: out <= 12'hee9;
      20'h0b669: out <= 12'hf87;
      20'h0b66a: out <= 12'hf87;
      20'h0b66b: out <= 12'hf87;
      20'h0b66c: out <= 12'hf87;
      20'h0b66d: out <= 12'hf87;
      20'h0b66e: out <= 12'hf87;
      20'h0b66f: out <= 12'hb27;
      20'h0b670: out <= 12'h000;
      20'h0b671: out <= 12'h000;
      20'h0b672: out <= 12'h000;
      20'h0b673: out <= 12'h000;
      20'h0b674: out <= 12'h000;
      20'h0b675: out <= 12'h000;
      20'h0b676: out <= 12'h000;
      20'h0b677: out <= 12'h000;
      20'h0b678: out <= 12'h777;
      20'h0b679: out <= 12'h555;
      20'h0b67a: out <= 12'h555;
      20'h0b67b: out <= 12'h555;
      20'h0b67c: out <= 12'h555;
      20'h0b67d: out <= 12'h555;
      20'h0b67e: out <= 12'h555;
      20'h0b67f: out <= 12'h555;
      20'h0b680: out <= 12'h555;
      20'h0b681: out <= 12'h555;
      20'h0b682: out <= 12'h555;
      20'h0b683: out <= 12'h555;
      20'h0b684: out <= 12'h555;
      20'h0b685: out <= 12'h555;
      20'h0b686: out <= 12'h555;
      20'h0b687: out <= 12'h777;
      20'h0b688: out <= 12'h000;
      20'h0b689: out <= 12'h000;
      20'h0b68a: out <= 12'h000;
      20'h0b68b: out <= 12'h000;
      20'h0b68c: out <= 12'h000;
      20'h0b68d: out <= 12'h000;
      20'h0b68e: out <= 12'h000;
      20'h0b68f: out <= 12'h000;
      20'h0b690: out <= 12'h000;
      20'h0b691: out <= 12'h000;
      20'h0b692: out <= 12'h000;
      20'h0b693: out <= 12'h000;
      20'h0b694: out <= 12'h000;
      20'h0b695: out <= 12'h000;
      20'h0b696: out <= 12'h000;
      20'h0b697: out <= 12'h000;
      20'h0b698: out <= 12'h000;
      20'h0b699: out <= 12'h000;
      20'h0b69a: out <= 12'h000;
      20'h0b69b: out <= 12'h000;
      20'h0b69c: out <= 12'h000;
      20'h0b69d: out <= 12'h000;
      20'h0b69e: out <= 12'h000;
      20'h0b69f: out <= 12'h000;
      20'h0b6a0: out <= 12'h000;
      20'h0b6a1: out <= 12'h000;
      20'h0b6a2: out <= 12'h000;
      20'h0b6a3: out <= 12'h000;
      20'h0b6a4: out <= 12'h000;
      20'h0b6a5: out <= 12'h000;
      20'h0b6a6: out <= 12'h000;
      20'h0b6a7: out <= 12'h000;
      20'h0b6a8: out <= 12'h088;
      20'h0b6a9: out <= 12'h088;
      20'h0b6aa: out <= 12'h088;
      20'h0b6ab: out <= 12'h088;
      20'h0b6ac: out <= 12'h088;
      20'h0b6ad: out <= 12'h088;
      20'h0b6ae: out <= 12'h088;
      20'h0b6af: out <= 12'h088;
      20'h0b6b0: out <= 12'h088;
      20'h0b6b1: out <= 12'h088;
      20'h0b6b2: out <= 12'h088;
      20'h0b6b3: out <= 12'h088;
      20'h0b6b4: out <= 12'h088;
      20'h0b6b5: out <= 12'h088;
      20'h0b6b6: out <= 12'h088;
      20'h0b6b7: out <= 12'h088;
      20'h0b6b8: out <= 12'h088;
      20'h0b6b9: out <= 12'h088;
      20'h0b6ba: out <= 12'h088;
      20'h0b6bb: out <= 12'h088;
      20'h0b6bc: out <= 12'h088;
      20'h0b6bd: out <= 12'h088;
      20'h0b6be: out <= 12'h088;
      20'h0b6bf: out <= 12'h088;
      20'h0b6c0: out <= 12'h088;
      20'h0b6c1: out <= 12'h088;
      20'h0b6c2: out <= 12'h088;
      20'h0b6c3: out <= 12'h088;
      20'h0b6c4: out <= 12'h088;
      20'h0b6c5: out <= 12'h088;
      20'h0b6c6: out <= 12'h088;
      20'h0b6c7: out <= 12'h088;
      20'h0b6c8: out <= 12'h088;
      20'h0b6c9: out <= 12'h088;
      20'h0b6ca: out <= 12'h088;
      20'h0b6cb: out <= 12'h088;
      20'h0b6cc: out <= 12'h088;
      20'h0b6cd: out <= 12'h088;
      20'h0b6ce: out <= 12'h088;
      20'h0b6cf: out <= 12'h088;
      20'h0b6d0: out <= 12'h088;
      20'h0b6d1: out <= 12'h088;
      20'h0b6d2: out <= 12'h088;
      20'h0b6d3: out <= 12'h088;
      20'h0b6d4: out <= 12'h088;
      20'h0b6d5: out <= 12'h088;
      20'h0b6d6: out <= 12'h088;
      20'h0b6d7: out <= 12'h088;
      20'h0b6d8: out <= 12'h088;
      20'h0b6d9: out <= 12'h088;
      20'h0b6da: out <= 12'h088;
      20'h0b6db: out <= 12'h088;
      20'h0b6dc: out <= 12'h088;
      20'h0b6dd: out <= 12'h088;
      20'h0b6de: out <= 12'h088;
      20'h0b6df: out <= 12'h088;
      20'h0b6e0: out <= 12'h088;
      20'h0b6e1: out <= 12'h088;
      20'h0b6e2: out <= 12'h088;
      20'h0b6e3: out <= 12'h088;
      20'h0b6e4: out <= 12'h088;
      20'h0b6e5: out <= 12'h088;
      20'h0b6e6: out <= 12'h088;
      20'h0b6e7: out <= 12'h088;
      20'h0b6e8: out <= 12'h088;
      20'h0b6e9: out <= 12'h088;
      20'h0b6ea: out <= 12'h088;
      20'h0b6eb: out <= 12'h088;
      20'h0b6ec: out <= 12'h088;
      20'h0b6ed: out <= 12'h088;
      20'h0b6ee: out <= 12'h088;
      20'h0b6ef: out <= 12'h088;
      20'h0b6f0: out <= 12'h088;
      20'h0b6f1: out <= 12'h088;
      20'h0b6f2: out <= 12'h088;
      20'h0b6f3: out <= 12'h088;
      20'h0b6f4: out <= 12'h088;
      20'h0b6f5: out <= 12'h088;
      20'h0b6f6: out <= 12'h088;
      20'h0b6f7: out <= 12'h088;
      20'h0b6f8: out <= 12'h088;
      20'h0b6f9: out <= 12'h088;
      20'h0b6fa: out <= 12'h088;
      20'h0b6fb: out <= 12'h088;
      20'h0b6fc: out <= 12'h088;
      20'h0b6fd: out <= 12'h088;
      20'h0b6fe: out <= 12'h088;
      20'h0b6ff: out <= 12'h088;
      20'h0b700: out <= 12'h088;
      20'h0b701: out <= 12'h088;
      20'h0b702: out <= 12'h088;
      20'h0b703: out <= 12'h088;
      20'h0b704: out <= 12'h088;
      20'h0b705: out <= 12'h088;
      20'h0b706: out <= 12'h088;
      20'h0b707: out <= 12'h088;
      20'h0b708: out <= 12'h088;
      20'h0b709: out <= 12'h088;
      20'h0b70a: out <= 12'h088;
      20'h0b70b: out <= 12'h088;
      20'h0b70c: out <= 12'h088;
      20'h0b70d: out <= 12'h088;
      20'h0b70e: out <= 12'h088;
      20'h0b70f: out <= 12'h088;
      20'h0b710: out <= 12'h088;
      20'h0b711: out <= 12'h222;
      20'h0b712: out <= 12'h222;
      20'h0b713: out <= 12'h222;
      20'h0b714: out <= 12'h222;
      20'h0b715: out <= 12'h222;
      20'h0b716: out <= 12'h222;
      20'h0b717: out <= 12'h222;
      20'h0b718: out <= 12'h222;
      20'h0b719: out <= 12'h222;
      20'h0b71a: out <= 12'h222;
      20'h0b71b: out <= 12'h222;
      20'h0b71c: out <= 12'hbb0;
      20'h0b71d: out <= 12'h222;
      20'h0b71e: out <= 12'h222;
      20'h0b71f: out <= 12'h222;
      20'h0b720: out <= 12'h222;
      20'h0b721: out <= 12'h222;
      20'h0b722: out <= 12'h222;
      20'h0b723: out <= 12'h222;
      20'h0b724: out <= 12'h222;
      20'h0b725: out <= 12'h222;
      20'h0b726: out <= 12'h222;
      20'h0b727: out <= 12'h222;
      20'h0b728: out <= 12'h603;
      20'h0b729: out <= 12'h603;
      20'h0b72a: out <= 12'h603;
      20'h0b72b: out <= 12'h603;
      20'h0b72c: out <= 12'h000;
      20'h0b72d: out <= 12'h000;
      20'h0b72e: out <= 12'h000;
      20'h0b72f: out <= 12'h000;
      20'h0b730: out <= 12'h000;
      20'h0b731: out <= 12'h000;
      20'h0b732: out <= 12'h000;
      20'h0b733: out <= 12'h000;
      20'h0b734: out <= 12'h000;
      20'h0b735: out <= 12'h000;
      20'h0b736: out <= 12'h000;
      20'h0b737: out <= 12'h000;
      20'h0b738: out <= 12'h000;
      20'h0b739: out <= 12'h000;
      20'h0b73a: out <= 12'h000;
      20'h0b73b: out <= 12'h000;
      20'h0b73c: out <= 12'h000;
      20'h0b73d: out <= 12'h000;
      20'h0b73e: out <= 12'h000;
      20'h0b73f: out <= 12'h000;
      20'h0b740: out <= 12'h000;
      20'h0b741: out <= 12'h000;
      20'h0b742: out <= 12'h000;
      20'h0b743: out <= 12'h000;
      20'h0b744: out <= 12'h000;
      20'h0b745: out <= 12'h000;
      20'h0b746: out <= 12'h000;
      20'h0b747: out <= 12'h000;
      20'h0b748: out <= 12'h000;
      20'h0b749: out <= 12'h000;
      20'h0b74a: out <= 12'h000;
      20'h0b74b: out <= 12'h000;
      20'h0b74c: out <= 12'h000;
      20'h0b74d: out <= 12'h000;
      20'h0b74e: out <= 12'h000;
      20'h0b74f: out <= 12'h000;
      20'h0b750: out <= 12'h000;
      20'h0b751: out <= 12'h000;
      20'h0b752: out <= 12'h000;
      20'h0b753: out <= 12'h000;
      20'h0b754: out <= 12'h000;
      20'h0b755: out <= 12'h000;
      20'h0b756: out <= 12'h000;
      20'h0b757: out <= 12'h000;
      20'h0b758: out <= 12'h000;
      20'h0b759: out <= 12'h000;
      20'h0b75a: out <= 12'h000;
      20'h0b75b: out <= 12'h000;
      20'h0b75c: out <= 12'h000;
      20'h0b75d: out <= 12'h000;
      20'h0b75e: out <= 12'h000;
      20'h0b75f: out <= 12'h000;
      20'h0b760: out <= 12'h000;
      20'h0b761: out <= 12'h000;
      20'h0b762: out <= 12'h000;
      20'h0b763: out <= 12'h000;
      20'h0b764: out <= 12'h000;
      20'h0b765: out <= 12'h000;
      20'h0b766: out <= 12'h000;
      20'h0b767: out <= 12'h000;
      20'h0b768: out <= 12'h000;
      20'h0b769: out <= 12'h000;
      20'h0b76a: out <= 12'h000;
      20'h0b76b: out <= 12'h000;
      20'h0b76c: out <= 12'h000;
      20'h0b76d: out <= 12'h000;
      20'h0b76e: out <= 12'h000;
      20'h0b76f: out <= 12'h000;
      20'h0b770: out <= 12'h000;
      20'h0b771: out <= 12'h000;
      20'h0b772: out <= 12'h000;
      20'h0b773: out <= 12'h000;
      20'h0b774: out <= 12'h000;
      20'h0b775: out <= 12'h000;
      20'h0b776: out <= 12'h000;
      20'h0b777: out <= 12'h000;
      20'h0b778: out <= 12'h000;
      20'h0b779: out <= 12'h000;
      20'h0b77a: out <= 12'h000;
      20'h0b77b: out <= 12'h000;
      20'h0b77c: out <= 12'h603;
      20'h0b77d: out <= 12'h603;
      20'h0b77e: out <= 12'h603;
      20'h0b77f: out <= 12'h603;
      20'h0b780: out <= 12'hb27;
      20'h0b781: out <= 12'hb27;
      20'h0b782: out <= 12'hb27;
      20'h0b783: out <= 12'hb27;
      20'h0b784: out <= 12'hb27;
      20'h0b785: out <= 12'hb27;
      20'h0b786: out <= 12'hb27;
      20'h0b787: out <= 12'hb27;
      20'h0b788: out <= 12'h000;
      20'h0b789: out <= 12'h000;
      20'h0b78a: out <= 12'h000;
      20'h0b78b: out <= 12'h000;
      20'h0b78c: out <= 12'h000;
      20'h0b78d: out <= 12'h000;
      20'h0b78e: out <= 12'h000;
      20'h0b78f: out <= 12'h000;
      20'h0b790: out <= 12'h777;
      20'h0b791: out <= 12'h555;
      20'h0b792: out <= 12'h555;
      20'h0b793: out <= 12'h555;
      20'h0b794: out <= 12'h555;
      20'h0b795: out <= 12'h555;
      20'h0b796: out <= 12'h555;
      20'h0b797: out <= 12'h555;
      20'h0b798: out <= 12'h555;
      20'h0b799: out <= 12'h555;
      20'h0b79a: out <= 12'h555;
      20'h0b79b: out <= 12'h555;
      20'h0b79c: out <= 12'h555;
      20'h0b79d: out <= 12'h555;
      20'h0b79e: out <= 12'h555;
      20'h0b79f: out <= 12'h777;
      20'h0b7a0: out <= 12'h000;
      20'h0b7a1: out <= 12'h000;
      20'h0b7a2: out <= 12'h000;
      20'h0b7a3: out <= 12'h000;
      20'h0b7a4: out <= 12'h000;
      20'h0b7a5: out <= 12'h000;
      20'h0b7a6: out <= 12'h000;
      20'h0b7a7: out <= 12'h000;
      20'h0b7a8: out <= 12'h000;
      20'h0b7a9: out <= 12'h000;
      20'h0b7aa: out <= 12'h000;
      20'h0b7ab: out <= 12'h000;
      20'h0b7ac: out <= 12'h000;
      20'h0b7ad: out <= 12'h000;
      20'h0b7ae: out <= 12'h000;
      20'h0b7af: out <= 12'h000;
      20'h0b7b0: out <= 12'h000;
      20'h0b7b1: out <= 12'h000;
      20'h0b7b2: out <= 12'h000;
      20'h0b7b3: out <= 12'h000;
      20'h0b7b4: out <= 12'h000;
      20'h0b7b5: out <= 12'h000;
      20'h0b7b6: out <= 12'h000;
      20'h0b7b7: out <= 12'h000;
      20'h0b7b8: out <= 12'h000;
      20'h0b7b9: out <= 12'h000;
      20'h0b7ba: out <= 12'h000;
      20'h0b7bb: out <= 12'h000;
      20'h0b7bc: out <= 12'h000;
      20'h0b7bd: out <= 12'h000;
      20'h0b7be: out <= 12'h000;
      20'h0b7bf: out <= 12'h000;
      20'h0b7c0: out <= 12'h088;
      20'h0b7c1: out <= 12'h088;
      20'h0b7c2: out <= 12'h088;
      20'h0b7c3: out <= 12'h088;
      20'h0b7c4: out <= 12'h088;
      20'h0b7c5: out <= 12'h088;
      20'h0b7c6: out <= 12'h088;
      20'h0b7c7: out <= 12'h088;
      20'h0b7c8: out <= 12'h088;
      20'h0b7c9: out <= 12'h088;
      20'h0b7ca: out <= 12'h088;
      20'h0b7cb: out <= 12'h088;
      20'h0b7cc: out <= 12'h088;
      20'h0b7cd: out <= 12'h088;
      20'h0b7ce: out <= 12'h088;
      20'h0b7cf: out <= 12'h088;
      20'h0b7d0: out <= 12'h088;
      20'h0b7d1: out <= 12'h088;
      20'h0b7d2: out <= 12'h088;
      20'h0b7d3: out <= 12'h088;
      20'h0b7d4: out <= 12'h088;
      20'h0b7d5: out <= 12'h088;
      20'h0b7d6: out <= 12'h088;
      20'h0b7d7: out <= 12'h088;
      20'h0b7d8: out <= 12'h088;
      20'h0b7d9: out <= 12'h088;
      20'h0b7da: out <= 12'h088;
      20'h0b7db: out <= 12'h088;
      20'h0b7dc: out <= 12'h088;
      20'h0b7dd: out <= 12'h088;
      20'h0b7de: out <= 12'h088;
      20'h0b7df: out <= 12'h088;
      20'h0b7e0: out <= 12'h088;
      20'h0b7e1: out <= 12'h088;
      20'h0b7e2: out <= 12'h088;
      20'h0b7e3: out <= 12'h088;
      20'h0b7e4: out <= 12'h088;
      20'h0b7e5: out <= 12'h088;
      20'h0b7e6: out <= 12'h088;
      20'h0b7e7: out <= 12'h088;
      20'h0b7e8: out <= 12'h088;
      20'h0b7e9: out <= 12'h088;
      20'h0b7ea: out <= 12'h088;
      20'h0b7eb: out <= 12'h088;
      20'h0b7ec: out <= 12'h088;
      20'h0b7ed: out <= 12'h088;
      20'h0b7ee: out <= 12'h088;
      20'h0b7ef: out <= 12'h088;
      20'h0b7f0: out <= 12'h088;
      20'h0b7f1: out <= 12'h088;
      20'h0b7f2: out <= 12'h088;
      20'h0b7f3: out <= 12'h088;
      20'h0b7f4: out <= 12'h088;
      20'h0b7f5: out <= 12'h088;
      20'h0b7f6: out <= 12'h088;
      20'h0b7f7: out <= 12'h088;
      20'h0b7f8: out <= 12'h088;
      20'h0b7f9: out <= 12'h088;
      20'h0b7fa: out <= 12'h088;
      20'h0b7fb: out <= 12'h088;
      20'h0b7fc: out <= 12'h088;
      20'h0b7fd: out <= 12'h088;
      20'h0b7fe: out <= 12'h088;
      20'h0b7ff: out <= 12'h088;
      20'h0b800: out <= 12'h088;
      20'h0b801: out <= 12'h088;
      20'h0b802: out <= 12'h088;
      20'h0b803: out <= 12'h088;
      20'h0b804: out <= 12'h088;
      20'h0b805: out <= 12'h088;
      20'h0b806: out <= 12'h088;
      20'h0b807: out <= 12'h088;
      20'h0b808: out <= 12'h088;
      20'h0b809: out <= 12'h088;
      20'h0b80a: out <= 12'h088;
      20'h0b80b: out <= 12'h088;
      20'h0b80c: out <= 12'h088;
      20'h0b80d: out <= 12'h088;
      20'h0b80e: out <= 12'h088;
      20'h0b80f: out <= 12'h088;
      20'h0b810: out <= 12'h088;
      20'h0b811: out <= 12'h088;
      20'h0b812: out <= 12'h088;
      20'h0b813: out <= 12'h088;
      20'h0b814: out <= 12'h088;
      20'h0b815: out <= 12'h088;
      20'h0b816: out <= 12'h088;
      20'h0b817: out <= 12'h088;
      20'h0b818: out <= 12'h088;
      20'h0b819: out <= 12'h088;
      20'h0b81a: out <= 12'h088;
      20'h0b81b: out <= 12'h088;
      20'h0b81c: out <= 12'h088;
      20'h0b81d: out <= 12'h088;
      20'h0b81e: out <= 12'h088;
      20'h0b81f: out <= 12'h088;
      20'h0b820: out <= 12'h088;
      20'h0b821: out <= 12'h088;
      20'h0b822: out <= 12'h088;
      20'h0b823: out <= 12'h088;
      20'h0b824: out <= 12'h088;
      20'h0b825: out <= 12'h088;
      20'h0b826: out <= 12'h088;
      20'h0b827: out <= 12'h088;
      20'h0b828: out <= 12'h088;
      20'h0b829: out <= 12'h222;
      20'h0b82a: out <= 12'h222;
      20'h0b82b: out <= 12'h222;
      20'h0b82c: out <= 12'h222;
      20'h0b82d: out <= 12'h222;
      20'h0b82e: out <= 12'h222;
      20'h0b82f: out <= 12'h222;
      20'h0b830: out <= 12'h222;
      20'h0b831: out <= 12'h222;
      20'h0b832: out <= 12'h222;
      20'h0b833: out <= 12'h660;
      20'h0b834: out <= 12'hee9;
      20'h0b835: out <= 12'h660;
      20'h0b836: out <= 12'h222;
      20'h0b837: out <= 12'h222;
      20'h0b838: out <= 12'h222;
      20'h0b839: out <= 12'h222;
      20'h0b83a: out <= 12'h222;
      20'h0b83b: out <= 12'h222;
      20'h0b83c: out <= 12'h222;
      20'h0b83d: out <= 12'h222;
      20'h0b83e: out <= 12'h222;
      20'h0b83f: out <= 12'h222;
      20'h0b840: out <= 12'h603;
      20'h0b841: out <= 12'h603;
      20'h0b842: out <= 12'h603;
      20'h0b843: out <= 12'h603;
      20'h0b844: out <= 12'h000;
      20'h0b845: out <= 12'hb27;
      20'h0b846: out <= 12'hb27;
      20'h0b847: out <= 12'hb27;
      20'h0b848: out <= 12'hb27;
      20'h0b849: out <= 12'hb27;
      20'h0b84a: out <= 12'h000;
      20'h0b84b: out <= 12'h000;
      20'h0b84c: out <= 12'h000;
      20'h0b84d: out <= 12'h000;
      20'h0b84e: out <= 12'h000;
      20'h0b84f: out <= 12'hb27;
      20'h0b850: out <= 12'hb27;
      20'h0b851: out <= 12'h000;
      20'h0b852: out <= 12'h000;
      20'h0b853: out <= 12'h000;
      20'h0b854: out <= 12'h000;
      20'h0b855: out <= 12'hb27;
      20'h0b856: out <= 12'hb27;
      20'h0b857: out <= 12'hb27;
      20'h0b858: out <= 12'hb27;
      20'h0b859: out <= 12'hb27;
      20'h0b85a: out <= 12'h000;
      20'h0b85b: out <= 12'h000;
      20'h0b85c: out <= 12'h000;
      20'h0b85d: out <= 12'hb27;
      20'h0b85e: out <= 12'hb27;
      20'h0b85f: out <= 12'hb27;
      20'h0b860: out <= 12'hb27;
      20'h0b861: out <= 12'hb27;
      20'h0b862: out <= 12'h000;
      20'h0b863: out <= 12'h000;
      20'h0b864: out <= 12'h000;
      20'h0b865: out <= 12'h000;
      20'h0b866: out <= 12'h000;
      20'h0b867: out <= 12'hb27;
      20'h0b868: out <= 12'hb27;
      20'h0b869: out <= 12'hb27;
      20'h0b86a: out <= 12'h000;
      20'h0b86b: out <= 12'h000;
      20'h0b86c: out <= 12'hb27;
      20'h0b86d: out <= 12'hb27;
      20'h0b86e: out <= 12'hb27;
      20'h0b86f: out <= 12'hb27;
      20'h0b870: out <= 12'hb27;
      20'h0b871: out <= 12'hb27;
      20'h0b872: out <= 12'hb27;
      20'h0b873: out <= 12'h000;
      20'h0b874: out <= 12'h000;
      20'h0b875: out <= 12'h000;
      20'h0b876: out <= 12'h000;
      20'h0b877: out <= 12'hb27;
      20'h0b878: out <= 12'hb27;
      20'h0b879: out <= 12'hb27;
      20'h0b87a: out <= 12'h000;
      20'h0b87b: out <= 12'h000;
      20'h0b87c: out <= 12'hb27;
      20'h0b87d: out <= 12'hb27;
      20'h0b87e: out <= 12'hb27;
      20'h0b87f: out <= 12'hb27;
      20'h0b880: out <= 12'hb27;
      20'h0b881: out <= 12'hb27;
      20'h0b882: out <= 12'hb27;
      20'h0b883: out <= 12'h000;
      20'h0b884: out <= 12'h000;
      20'h0b885: out <= 12'hb27;
      20'h0b886: out <= 12'hb27;
      20'h0b887: out <= 12'hb27;
      20'h0b888: out <= 12'hb27;
      20'h0b889: out <= 12'hb27;
      20'h0b88a: out <= 12'h000;
      20'h0b88b: out <= 12'h000;
      20'h0b88c: out <= 12'h000;
      20'h0b88d: out <= 12'hb27;
      20'h0b88e: out <= 12'hb27;
      20'h0b88f: out <= 12'hb27;
      20'h0b890: out <= 12'hb27;
      20'h0b891: out <= 12'hb27;
      20'h0b892: out <= 12'h000;
      20'h0b893: out <= 12'h000;
      20'h0b894: out <= 12'h603;
      20'h0b895: out <= 12'h603;
      20'h0b896: out <= 12'h603;
      20'h0b897: out <= 12'h603;
      20'h0b898: out <= 12'hee9;
      20'h0b899: out <= 12'hee9;
      20'h0b89a: out <= 12'hee9;
      20'h0b89b: out <= 12'hee9;
      20'h0b89c: out <= 12'hee9;
      20'h0b89d: out <= 12'hee9;
      20'h0b89e: out <= 12'hee9;
      20'h0b89f: out <= 12'hb27;
      20'h0b8a0: out <= 12'h000;
      20'h0b8a1: out <= 12'h000;
      20'h0b8a2: out <= 12'h000;
      20'h0b8a3: out <= 12'h000;
      20'h0b8a4: out <= 12'h000;
      20'h0b8a5: out <= 12'h000;
      20'h0b8a6: out <= 12'h000;
      20'h0b8a7: out <= 12'h000;
      20'h0b8a8: out <= 12'h777;
      20'h0b8a9: out <= 12'h555;
      20'h0b8aa: out <= 12'h555;
      20'h0b8ab: out <= 12'h555;
      20'h0b8ac: out <= 12'h555;
      20'h0b8ad: out <= 12'h555;
      20'h0b8ae: out <= 12'h555;
      20'h0b8af: out <= 12'h555;
      20'h0b8b0: out <= 12'h555;
      20'h0b8b1: out <= 12'h555;
      20'h0b8b2: out <= 12'h555;
      20'h0b8b3: out <= 12'h555;
      20'h0b8b4: out <= 12'h555;
      20'h0b8b5: out <= 12'h555;
      20'h0b8b6: out <= 12'h555;
      20'h0b8b7: out <= 12'h777;
      20'h0b8b8: out <= 12'h000;
      20'h0b8b9: out <= 12'h000;
      20'h0b8ba: out <= 12'h000;
      20'h0b8bb: out <= 12'h000;
      20'h0b8bc: out <= 12'h000;
      20'h0b8bd: out <= 12'h000;
      20'h0b8be: out <= 12'h000;
      20'h0b8bf: out <= 12'h000;
      20'h0b8c0: out <= 12'hfa9;
      20'h0b8c1: out <= 12'hfa9;
      20'h0b8c2: out <= 12'hfa9;
      20'h0b8c3: out <= 12'hfa9;
      20'h0b8c4: out <= 12'hfa9;
      20'h0b8c5: out <= 12'hfa9;
      20'h0b8c6: out <= 12'hfa9;
      20'h0b8c7: out <= 12'hfa9;
      20'h0b8c8: out <= 12'hf76;
      20'h0b8c9: out <= 12'hf76;
      20'h0b8ca: out <= 12'hf76;
      20'h0b8cb: out <= 12'hf76;
      20'h0b8cc: out <= 12'hf76;
      20'h0b8cd: out <= 12'hf76;
      20'h0b8ce: out <= 12'hf76;
      20'h0b8cf: out <= 12'hf76;
      20'h0b8d0: out <= 12'h000;
      20'h0b8d1: out <= 12'h000;
      20'h0b8d2: out <= 12'h000;
      20'h0b8d3: out <= 12'h000;
      20'h0b8d4: out <= 12'h000;
      20'h0b8d5: out <= 12'h000;
      20'h0b8d6: out <= 12'h000;
      20'h0b8d7: out <= 12'h000;
      20'h0b8d8: out <= 12'h088;
      20'h0b8d9: out <= 12'h088;
      20'h0b8da: out <= 12'h088;
      20'h0b8db: out <= 12'h088;
      20'h0b8dc: out <= 12'h088;
      20'h0b8dd: out <= 12'h088;
      20'h0b8de: out <= 12'h088;
      20'h0b8df: out <= 12'h088;
      20'h0b8e0: out <= 12'h088;
      20'h0b8e1: out <= 12'h088;
      20'h0b8e2: out <= 12'h088;
      20'h0b8e3: out <= 12'h088;
      20'h0b8e4: out <= 12'h088;
      20'h0b8e5: out <= 12'h088;
      20'h0b8e6: out <= 12'h088;
      20'h0b8e7: out <= 12'h088;
      20'h0b8e8: out <= 12'h088;
      20'h0b8e9: out <= 12'h088;
      20'h0b8ea: out <= 12'h088;
      20'h0b8eb: out <= 12'h088;
      20'h0b8ec: out <= 12'h088;
      20'h0b8ed: out <= 12'h088;
      20'h0b8ee: out <= 12'h088;
      20'h0b8ef: out <= 12'h088;
      20'h0b8f0: out <= 12'h088;
      20'h0b8f1: out <= 12'h088;
      20'h0b8f2: out <= 12'h088;
      20'h0b8f3: out <= 12'h088;
      20'h0b8f4: out <= 12'h088;
      20'h0b8f5: out <= 12'h088;
      20'h0b8f6: out <= 12'h088;
      20'h0b8f7: out <= 12'h088;
      20'h0b8f8: out <= 12'h088;
      20'h0b8f9: out <= 12'h088;
      20'h0b8fa: out <= 12'h088;
      20'h0b8fb: out <= 12'h088;
      20'h0b8fc: out <= 12'h088;
      20'h0b8fd: out <= 12'h088;
      20'h0b8fe: out <= 12'h088;
      20'h0b8ff: out <= 12'h088;
      20'h0b900: out <= 12'h088;
      20'h0b901: out <= 12'h088;
      20'h0b902: out <= 12'h088;
      20'h0b903: out <= 12'h088;
      20'h0b904: out <= 12'h088;
      20'h0b905: out <= 12'h088;
      20'h0b906: out <= 12'h088;
      20'h0b907: out <= 12'h088;
      20'h0b908: out <= 12'h088;
      20'h0b909: out <= 12'h088;
      20'h0b90a: out <= 12'h088;
      20'h0b90b: out <= 12'h088;
      20'h0b90c: out <= 12'h088;
      20'h0b90d: out <= 12'h088;
      20'h0b90e: out <= 12'h088;
      20'h0b90f: out <= 12'h088;
      20'h0b910: out <= 12'h088;
      20'h0b911: out <= 12'h088;
      20'h0b912: out <= 12'h088;
      20'h0b913: out <= 12'h088;
      20'h0b914: out <= 12'h088;
      20'h0b915: out <= 12'h088;
      20'h0b916: out <= 12'h088;
      20'h0b917: out <= 12'h088;
      20'h0b918: out <= 12'h088;
      20'h0b919: out <= 12'h088;
      20'h0b91a: out <= 12'h088;
      20'h0b91b: out <= 12'h088;
      20'h0b91c: out <= 12'h088;
      20'h0b91d: out <= 12'h088;
      20'h0b91e: out <= 12'h088;
      20'h0b91f: out <= 12'h088;
      20'h0b920: out <= 12'h088;
      20'h0b921: out <= 12'h088;
      20'h0b922: out <= 12'h088;
      20'h0b923: out <= 12'h088;
      20'h0b924: out <= 12'h088;
      20'h0b925: out <= 12'h088;
      20'h0b926: out <= 12'h088;
      20'h0b927: out <= 12'h088;
      20'h0b928: out <= 12'h088;
      20'h0b929: out <= 12'h088;
      20'h0b92a: out <= 12'h088;
      20'h0b92b: out <= 12'h088;
      20'h0b92c: out <= 12'h088;
      20'h0b92d: out <= 12'h088;
      20'h0b92e: out <= 12'h088;
      20'h0b92f: out <= 12'h088;
      20'h0b930: out <= 12'h088;
      20'h0b931: out <= 12'h088;
      20'h0b932: out <= 12'h088;
      20'h0b933: out <= 12'h088;
      20'h0b934: out <= 12'h088;
      20'h0b935: out <= 12'h088;
      20'h0b936: out <= 12'h088;
      20'h0b937: out <= 12'h088;
      20'h0b938: out <= 12'h088;
      20'h0b939: out <= 12'h088;
      20'h0b93a: out <= 12'h088;
      20'h0b93b: out <= 12'h088;
      20'h0b93c: out <= 12'h088;
      20'h0b93d: out <= 12'h088;
      20'h0b93e: out <= 12'h088;
      20'h0b93f: out <= 12'h088;
      20'h0b940: out <= 12'h088;
      20'h0b941: out <= 12'h222;
      20'h0b942: out <= 12'h222;
      20'h0b943: out <= 12'h222;
      20'h0b944: out <= 12'h222;
      20'h0b945: out <= 12'h222;
      20'h0b946: out <= 12'h222;
      20'h0b947: out <= 12'h222;
      20'h0b948: out <= 12'h222;
      20'h0b949: out <= 12'h222;
      20'h0b94a: out <= 12'h660;
      20'h0b94b: out <= 12'hbb0;
      20'h0b94c: out <= 12'hee9;
      20'h0b94d: out <= 12'hbb0;
      20'h0b94e: out <= 12'h660;
      20'h0b94f: out <= 12'h222;
      20'h0b950: out <= 12'h222;
      20'h0b951: out <= 12'h222;
      20'h0b952: out <= 12'h222;
      20'h0b953: out <= 12'h222;
      20'h0b954: out <= 12'h222;
      20'h0b955: out <= 12'h222;
      20'h0b956: out <= 12'h222;
      20'h0b957: out <= 12'h222;
      20'h0b958: out <= 12'h603;
      20'h0b959: out <= 12'h603;
      20'h0b95a: out <= 12'h603;
      20'h0b95b: out <= 12'h603;
      20'h0b95c: out <= 12'hb27;
      20'h0b95d: out <= 12'hb27;
      20'h0b95e: out <= 12'hb27;
      20'h0b95f: out <= 12'hb27;
      20'h0b960: out <= 12'hb27;
      20'h0b961: out <= 12'hb27;
      20'h0b962: out <= 12'hb27;
      20'h0b963: out <= 12'h000;
      20'h0b964: out <= 12'h000;
      20'h0b965: out <= 12'h000;
      20'h0b966: out <= 12'h000;
      20'h0b967: out <= 12'hb27;
      20'h0b968: out <= 12'hb27;
      20'h0b969: out <= 12'h000;
      20'h0b96a: out <= 12'h000;
      20'h0b96b: out <= 12'h000;
      20'h0b96c: out <= 12'hb27;
      20'h0b96d: out <= 12'hb27;
      20'h0b96e: out <= 12'hb27;
      20'h0b96f: out <= 12'hb27;
      20'h0b970: out <= 12'hb27;
      20'h0b971: out <= 12'hb27;
      20'h0b972: out <= 12'hb27;
      20'h0b973: out <= 12'h000;
      20'h0b974: out <= 12'hb27;
      20'h0b975: out <= 12'hb27;
      20'h0b976: out <= 12'hb27;
      20'h0b977: out <= 12'hb27;
      20'h0b978: out <= 12'hb27;
      20'h0b979: out <= 12'hb27;
      20'h0b97a: out <= 12'hb27;
      20'h0b97b: out <= 12'h000;
      20'h0b97c: out <= 12'h000;
      20'h0b97d: out <= 12'h000;
      20'h0b97e: out <= 12'h000;
      20'h0b97f: out <= 12'hb27;
      20'h0b980: out <= 12'hb27;
      20'h0b981: out <= 12'hb27;
      20'h0b982: out <= 12'h000;
      20'h0b983: out <= 12'h000;
      20'h0b984: out <= 12'hb27;
      20'h0b985: out <= 12'hb27;
      20'h0b986: out <= 12'hb27;
      20'h0b987: out <= 12'hb27;
      20'h0b988: out <= 12'hb27;
      20'h0b989: out <= 12'hb27;
      20'h0b98a: out <= 12'hb27;
      20'h0b98b: out <= 12'h000;
      20'h0b98c: out <= 12'h000;
      20'h0b98d: out <= 12'h000;
      20'h0b98e: out <= 12'hb27;
      20'h0b98f: out <= 12'hb27;
      20'h0b990: out <= 12'hb27;
      20'h0b991: out <= 12'hb27;
      20'h0b992: out <= 12'h000;
      20'h0b993: out <= 12'h000;
      20'h0b994: out <= 12'hb27;
      20'h0b995: out <= 12'hb27;
      20'h0b996: out <= 12'hb27;
      20'h0b997: out <= 12'hb27;
      20'h0b998: out <= 12'hb27;
      20'h0b999: out <= 12'hb27;
      20'h0b99a: out <= 12'hb27;
      20'h0b99b: out <= 12'h000;
      20'h0b99c: out <= 12'hb27;
      20'h0b99d: out <= 12'hb27;
      20'h0b99e: out <= 12'hb27;
      20'h0b99f: out <= 12'hb27;
      20'h0b9a0: out <= 12'hb27;
      20'h0b9a1: out <= 12'hb27;
      20'h0b9a2: out <= 12'hb27;
      20'h0b9a3: out <= 12'h000;
      20'h0b9a4: out <= 12'hb27;
      20'h0b9a5: out <= 12'hb27;
      20'h0b9a6: out <= 12'hb27;
      20'h0b9a7: out <= 12'hb27;
      20'h0b9a8: out <= 12'hb27;
      20'h0b9a9: out <= 12'hb27;
      20'h0b9aa: out <= 12'hb27;
      20'h0b9ab: out <= 12'h000;
      20'h0b9ac: out <= 12'h603;
      20'h0b9ad: out <= 12'h603;
      20'h0b9ae: out <= 12'h603;
      20'h0b9af: out <= 12'h603;
      20'h0b9b0: out <= 12'hee9;
      20'h0b9b1: out <= 12'hf87;
      20'h0b9b2: out <= 12'hf87;
      20'h0b9b3: out <= 12'hf87;
      20'h0b9b4: out <= 12'hf87;
      20'h0b9b5: out <= 12'hf87;
      20'h0b9b6: out <= 12'hf87;
      20'h0b9b7: out <= 12'hb27;
      20'h0b9b8: out <= 12'h000;
      20'h0b9b9: out <= 12'h000;
      20'h0b9ba: out <= 12'h000;
      20'h0b9bb: out <= 12'h000;
      20'h0b9bc: out <= 12'h000;
      20'h0b9bd: out <= 12'h000;
      20'h0b9be: out <= 12'h000;
      20'h0b9bf: out <= 12'h000;
      20'h0b9c0: out <= 12'h777;
      20'h0b9c1: out <= 12'h555;
      20'h0b9c2: out <= 12'h555;
      20'h0b9c3: out <= 12'h555;
      20'h0b9c4: out <= 12'h555;
      20'h0b9c5: out <= 12'h555;
      20'h0b9c6: out <= 12'h555;
      20'h0b9c7: out <= 12'h555;
      20'h0b9c8: out <= 12'h555;
      20'h0b9c9: out <= 12'h555;
      20'h0b9ca: out <= 12'h555;
      20'h0b9cb: out <= 12'h555;
      20'h0b9cc: out <= 12'h555;
      20'h0b9cd: out <= 12'h555;
      20'h0b9ce: out <= 12'h555;
      20'h0b9cf: out <= 12'h777;
      20'h0b9d0: out <= 12'h000;
      20'h0b9d1: out <= 12'h000;
      20'h0b9d2: out <= 12'hf87;
      20'h0b9d3: out <= 12'h000;
      20'h0b9d4: out <= 12'h000;
      20'h0b9d5: out <= 12'h000;
      20'h0b9d6: out <= 12'hf87;
      20'h0b9d7: out <= 12'h000;
      20'h0b9d8: out <= 12'hfa9;
      20'h0b9d9: out <= 12'hfa9;
      20'h0b9da: out <= 12'hfa9;
      20'h0b9db: out <= 12'hfa9;
      20'h0b9dc: out <= 12'hfa9;
      20'h0b9dd: out <= 12'hfa9;
      20'h0b9de: out <= 12'hfa9;
      20'h0b9df: out <= 12'hfa9;
      20'h0b9e0: out <= 12'hf76;
      20'h0b9e1: out <= 12'hf76;
      20'h0b9e2: out <= 12'hf76;
      20'h0b9e3: out <= 12'hf76;
      20'h0b9e4: out <= 12'hf76;
      20'h0b9e5: out <= 12'hf76;
      20'h0b9e6: out <= 12'hf76;
      20'h0b9e7: out <= 12'hf76;
      20'h0b9e8: out <= 12'h000;
      20'h0b9e9: out <= 12'h000;
      20'h0b9ea: out <= 12'h000;
      20'h0b9eb: out <= 12'h000;
      20'h0b9ec: out <= 12'h000;
      20'h0b9ed: out <= 12'h000;
      20'h0b9ee: out <= 12'h000;
      20'h0b9ef: out <= 12'h000;
      20'h0b9f0: out <= 12'h088;
      20'h0b9f1: out <= 12'h088;
      20'h0b9f2: out <= 12'h088;
      20'h0b9f3: out <= 12'h088;
      20'h0b9f4: out <= 12'h088;
      20'h0b9f5: out <= 12'h088;
      20'h0b9f6: out <= 12'h088;
      20'h0b9f7: out <= 12'h088;
      20'h0b9f8: out <= 12'h088;
      20'h0b9f9: out <= 12'h088;
      20'h0b9fa: out <= 12'h088;
      20'h0b9fb: out <= 12'h088;
      20'h0b9fc: out <= 12'h088;
      20'h0b9fd: out <= 12'h088;
      20'h0b9fe: out <= 12'h088;
      20'h0b9ff: out <= 12'h088;
      20'h0ba00: out <= 12'h088;
      20'h0ba01: out <= 12'h088;
      20'h0ba02: out <= 12'h088;
      20'h0ba03: out <= 12'h088;
      20'h0ba04: out <= 12'h088;
      20'h0ba05: out <= 12'h088;
      20'h0ba06: out <= 12'h088;
      20'h0ba07: out <= 12'h088;
      20'h0ba08: out <= 12'h088;
      20'h0ba09: out <= 12'h088;
      20'h0ba0a: out <= 12'h088;
      20'h0ba0b: out <= 12'h088;
      20'h0ba0c: out <= 12'h088;
      20'h0ba0d: out <= 12'h088;
      20'h0ba0e: out <= 12'h088;
      20'h0ba0f: out <= 12'h088;
      20'h0ba10: out <= 12'h088;
      20'h0ba11: out <= 12'h088;
      20'h0ba12: out <= 12'h088;
      20'h0ba13: out <= 12'h088;
      20'h0ba14: out <= 12'h088;
      20'h0ba15: out <= 12'h088;
      20'h0ba16: out <= 12'h088;
      20'h0ba17: out <= 12'h088;
      20'h0ba18: out <= 12'h088;
      20'h0ba19: out <= 12'h088;
      20'h0ba1a: out <= 12'h088;
      20'h0ba1b: out <= 12'h088;
      20'h0ba1c: out <= 12'h088;
      20'h0ba1d: out <= 12'h088;
      20'h0ba1e: out <= 12'h088;
      20'h0ba1f: out <= 12'h088;
      20'h0ba20: out <= 12'h088;
      20'h0ba21: out <= 12'h088;
      20'h0ba22: out <= 12'h088;
      20'h0ba23: out <= 12'h088;
      20'h0ba24: out <= 12'h088;
      20'h0ba25: out <= 12'h088;
      20'h0ba26: out <= 12'h088;
      20'h0ba27: out <= 12'h088;
      20'h0ba28: out <= 12'h088;
      20'h0ba29: out <= 12'h088;
      20'h0ba2a: out <= 12'h088;
      20'h0ba2b: out <= 12'h088;
      20'h0ba2c: out <= 12'h088;
      20'h0ba2d: out <= 12'h088;
      20'h0ba2e: out <= 12'h088;
      20'h0ba2f: out <= 12'h088;
      20'h0ba30: out <= 12'h088;
      20'h0ba31: out <= 12'h088;
      20'h0ba32: out <= 12'h088;
      20'h0ba33: out <= 12'h088;
      20'h0ba34: out <= 12'h088;
      20'h0ba35: out <= 12'h088;
      20'h0ba36: out <= 12'h088;
      20'h0ba37: out <= 12'h088;
      20'h0ba38: out <= 12'h088;
      20'h0ba39: out <= 12'h088;
      20'h0ba3a: out <= 12'h088;
      20'h0ba3b: out <= 12'h088;
      20'h0ba3c: out <= 12'h088;
      20'h0ba3d: out <= 12'h088;
      20'h0ba3e: out <= 12'h088;
      20'h0ba3f: out <= 12'h088;
      20'h0ba40: out <= 12'h088;
      20'h0ba41: out <= 12'h088;
      20'h0ba42: out <= 12'h088;
      20'h0ba43: out <= 12'h088;
      20'h0ba44: out <= 12'h088;
      20'h0ba45: out <= 12'h088;
      20'h0ba46: out <= 12'h088;
      20'h0ba47: out <= 12'h088;
      20'h0ba48: out <= 12'h088;
      20'h0ba49: out <= 12'h088;
      20'h0ba4a: out <= 12'h088;
      20'h0ba4b: out <= 12'h088;
      20'h0ba4c: out <= 12'h088;
      20'h0ba4d: out <= 12'h088;
      20'h0ba4e: out <= 12'h088;
      20'h0ba4f: out <= 12'h088;
      20'h0ba50: out <= 12'h088;
      20'h0ba51: out <= 12'h088;
      20'h0ba52: out <= 12'h088;
      20'h0ba53: out <= 12'h088;
      20'h0ba54: out <= 12'h088;
      20'h0ba55: out <= 12'h088;
      20'h0ba56: out <= 12'h088;
      20'h0ba57: out <= 12'h088;
      20'h0ba58: out <= 12'h088;
      20'h0ba59: out <= 12'h222;
      20'h0ba5a: out <= 12'h222;
      20'h0ba5b: out <= 12'h222;
      20'h0ba5c: out <= 12'h222;
      20'h0ba5d: out <= 12'h222;
      20'h0ba5e: out <= 12'h222;
      20'h0ba5f: out <= 12'h222;
      20'h0ba60: out <= 12'h222;
      20'h0ba61: out <= 12'h660;
      20'h0ba62: out <= 12'hbb0;
      20'h0ba63: out <= 12'hee9;
      20'h0ba64: out <= 12'hee9;
      20'h0ba65: out <= 12'hee9;
      20'h0ba66: out <= 12'hbb0;
      20'h0ba67: out <= 12'h660;
      20'h0ba68: out <= 12'h222;
      20'h0ba69: out <= 12'h222;
      20'h0ba6a: out <= 12'h222;
      20'h0ba6b: out <= 12'h222;
      20'h0ba6c: out <= 12'h222;
      20'h0ba6d: out <= 12'h222;
      20'h0ba6e: out <= 12'h222;
      20'h0ba6f: out <= 12'h222;
      20'h0ba70: out <= 12'h603;
      20'h0ba71: out <= 12'h603;
      20'h0ba72: out <= 12'h603;
      20'h0ba73: out <= 12'h603;
      20'h0ba74: out <= 12'hf87;
      20'h0ba75: out <= 12'hf87;
      20'h0ba76: out <= 12'h000;
      20'h0ba77: out <= 12'h000;
      20'h0ba78: out <= 12'h000;
      20'h0ba79: out <= 12'hf87;
      20'h0ba7a: out <= 12'hf87;
      20'h0ba7b: out <= 12'h000;
      20'h0ba7c: out <= 12'h000;
      20'h0ba7d: out <= 12'h000;
      20'h0ba7e: out <= 12'hf87;
      20'h0ba7f: out <= 12'hf87;
      20'h0ba80: out <= 12'hf87;
      20'h0ba81: out <= 12'h000;
      20'h0ba82: out <= 12'h000;
      20'h0ba83: out <= 12'h000;
      20'h0ba84: out <= 12'hf87;
      20'h0ba85: out <= 12'hf87;
      20'h0ba86: out <= 12'h000;
      20'h0ba87: out <= 12'h000;
      20'h0ba88: out <= 12'h000;
      20'h0ba89: out <= 12'hf87;
      20'h0ba8a: out <= 12'hf87;
      20'h0ba8b: out <= 12'h000;
      20'h0ba8c: out <= 12'hf87;
      20'h0ba8d: out <= 12'hf87;
      20'h0ba8e: out <= 12'h000;
      20'h0ba8f: out <= 12'h000;
      20'h0ba90: out <= 12'h000;
      20'h0ba91: out <= 12'hf87;
      20'h0ba92: out <= 12'hf87;
      20'h0ba93: out <= 12'h000;
      20'h0ba94: out <= 12'h000;
      20'h0ba95: out <= 12'h000;
      20'h0ba96: out <= 12'hf87;
      20'h0ba97: out <= 12'hf87;
      20'h0ba98: out <= 12'hf87;
      20'h0ba99: out <= 12'hf87;
      20'h0ba9a: out <= 12'h000;
      20'h0ba9b: out <= 12'h000;
      20'h0ba9c: out <= 12'hf87;
      20'h0ba9d: out <= 12'hf87;
      20'h0ba9e: out <= 12'h000;
      20'h0ba9f: out <= 12'h000;
      20'h0baa0: out <= 12'h000;
      20'h0baa1: out <= 12'h000;
      20'h0baa2: out <= 12'h000;
      20'h0baa3: out <= 12'h000;
      20'h0baa4: out <= 12'h000;
      20'h0baa5: out <= 12'hf87;
      20'h0baa6: out <= 12'hf87;
      20'h0baa7: out <= 12'hf87;
      20'h0baa8: out <= 12'h000;
      20'h0baa9: out <= 12'h000;
      20'h0baaa: out <= 12'h000;
      20'h0baab: out <= 12'h000;
      20'h0baac: out <= 12'hf87;
      20'h0baad: out <= 12'hf87;
      20'h0baae: out <= 12'h000;
      20'h0baaf: out <= 12'h000;
      20'h0bab0: out <= 12'h000;
      20'h0bab1: out <= 12'hf87;
      20'h0bab2: out <= 12'hf87;
      20'h0bab3: out <= 12'h000;
      20'h0bab4: out <= 12'hf87;
      20'h0bab5: out <= 12'hf87;
      20'h0bab6: out <= 12'h000;
      20'h0bab7: out <= 12'h000;
      20'h0bab8: out <= 12'h000;
      20'h0bab9: out <= 12'hf87;
      20'h0baba: out <= 12'hf87;
      20'h0babb: out <= 12'h000;
      20'h0babc: out <= 12'hf87;
      20'h0babd: out <= 12'hf87;
      20'h0babe: out <= 12'h000;
      20'h0babf: out <= 12'h000;
      20'h0bac0: out <= 12'h000;
      20'h0bac1: out <= 12'hf87;
      20'h0bac2: out <= 12'hf87;
      20'h0bac3: out <= 12'h000;
      20'h0bac4: out <= 12'h603;
      20'h0bac5: out <= 12'h603;
      20'h0bac6: out <= 12'h603;
      20'h0bac7: out <= 12'h603;
      20'h0bac8: out <= 12'hee9;
      20'h0bac9: out <= 12'hf87;
      20'h0baca: out <= 12'hee9;
      20'h0bacb: out <= 12'hee9;
      20'h0bacc: out <= 12'hee9;
      20'h0bacd: out <= 12'hb27;
      20'h0bace: out <= 12'hf87;
      20'h0bacf: out <= 12'hb27;
      20'h0bad0: out <= 12'h000;
      20'h0bad1: out <= 12'h000;
      20'h0bad2: out <= 12'h000;
      20'h0bad3: out <= 12'h000;
      20'h0bad4: out <= 12'h000;
      20'h0bad5: out <= 12'h000;
      20'h0bad6: out <= 12'h000;
      20'h0bad7: out <= 12'h000;
      20'h0bad8: out <= 12'h777;
      20'h0bad9: out <= 12'h555;
      20'h0bada: out <= 12'h555;
      20'h0badb: out <= 12'h555;
      20'h0badc: out <= 12'h555;
      20'h0badd: out <= 12'h555;
      20'h0bade: out <= 12'h555;
      20'h0badf: out <= 12'h555;
      20'h0bae0: out <= 12'h555;
      20'h0bae1: out <= 12'h555;
      20'h0bae2: out <= 12'h555;
      20'h0bae3: out <= 12'h555;
      20'h0bae4: out <= 12'h555;
      20'h0bae5: out <= 12'h555;
      20'h0bae6: out <= 12'h555;
      20'h0bae7: out <= 12'h777;
      20'h0bae8: out <= 12'h000;
      20'h0bae9: out <= 12'h000;
      20'h0baea: out <= 12'h000;
      20'h0baeb: out <= 12'hf87;
      20'h0baec: out <= 12'h000;
      20'h0baed: out <= 12'hf87;
      20'h0baee: out <= 12'h000;
      20'h0baef: out <= 12'h000;
      20'h0baf0: out <= 12'hfa9;
      20'h0baf1: out <= 12'hfa9;
      20'h0baf2: out <= 12'hfa9;
      20'h0baf3: out <= 12'hfa9;
      20'h0baf4: out <= 12'hfa9;
      20'h0baf5: out <= 12'hfa9;
      20'h0baf6: out <= 12'hfa9;
      20'h0baf7: out <= 12'hfa9;
      20'h0baf8: out <= 12'hf76;
      20'h0baf9: out <= 12'hf76;
      20'h0bafa: out <= 12'hf76;
      20'h0bafb: out <= 12'hf76;
      20'h0bafc: out <= 12'hf76;
      20'h0bafd: out <= 12'hf76;
      20'h0bafe: out <= 12'hf76;
      20'h0baff: out <= 12'hf76;
      20'h0bb00: out <= 12'h000;
      20'h0bb01: out <= 12'h000;
      20'h0bb02: out <= 12'h000;
      20'h0bb03: out <= 12'h000;
      20'h0bb04: out <= 12'h000;
      20'h0bb05: out <= 12'h000;
      20'h0bb06: out <= 12'h000;
      20'h0bb07: out <= 12'h000;
      20'h0bb08: out <= 12'h088;
      20'h0bb09: out <= 12'h088;
      20'h0bb0a: out <= 12'h088;
      20'h0bb0b: out <= 12'h088;
      20'h0bb0c: out <= 12'h088;
      20'h0bb0d: out <= 12'h088;
      20'h0bb0e: out <= 12'h088;
      20'h0bb0f: out <= 12'h088;
      20'h0bb10: out <= 12'h088;
      20'h0bb11: out <= 12'h088;
      20'h0bb12: out <= 12'h088;
      20'h0bb13: out <= 12'h088;
      20'h0bb14: out <= 12'h088;
      20'h0bb15: out <= 12'h088;
      20'h0bb16: out <= 12'h088;
      20'h0bb17: out <= 12'h088;
      20'h0bb18: out <= 12'h088;
      20'h0bb19: out <= 12'h088;
      20'h0bb1a: out <= 12'h088;
      20'h0bb1b: out <= 12'h088;
      20'h0bb1c: out <= 12'h088;
      20'h0bb1d: out <= 12'h088;
      20'h0bb1e: out <= 12'h088;
      20'h0bb1f: out <= 12'h088;
      20'h0bb20: out <= 12'h088;
      20'h0bb21: out <= 12'h088;
      20'h0bb22: out <= 12'h088;
      20'h0bb23: out <= 12'h088;
      20'h0bb24: out <= 12'h088;
      20'h0bb25: out <= 12'h088;
      20'h0bb26: out <= 12'h088;
      20'h0bb27: out <= 12'h088;
      20'h0bb28: out <= 12'h088;
      20'h0bb29: out <= 12'h088;
      20'h0bb2a: out <= 12'h088;
      20'h0bb2b: out <= 12'h088;
      20'h0bb2c: out <= 12'h088;
      20'h0bb2d: out <= 12'h088;
      20'h0bb2e: out <= 12'h088;
      20'h0bb2f: out <= 12'h088;
      20'h0bb30: out <= 12'h088;
      20'h0bb31: out <= 12'h088;
      20'h0bb32: out <= 12'h088;
      20'h0bb33: out <= 12'h088;
      20'h0bb34: out <= 12'h088;
      20'h0bb35: out <= 12'h088;
      20'h0bb36: out <= 12'h088;
      20'h0bb37: out <= 12'h088;
      20'h0bb38: out <= 12'h088;
      20'h0bb39: out <= 12'h088;
      20'h0bb3a: out <= 12'h088;
      20'h0bb3b: out <= 12'h088;
      20'h0bb3c: out <= 12'h088;
      20'h0bb3d: out <= 12'h088;
      20'h0bb3e: out <= 12'h088;
      20'h0bb3f: out <= 12'h088;
      20'h0bb40: out <= 12'h088;
      20'h0bb41: out <= 12'h088;
      20'h0bb42: out <= 12'h088;
      20'h0bb43: out <= 12'h088;
      20'h0bb44: out <= 12'h088;
      20'h0bb45: out <= 12'h088;
      20'h0bb46: out <= 12'h088;
      20'h0bb47: out <= 12'h088;
      20'h0bb48: out <= 12'h088;
      20'h0bb49: out <= 12'h088;
      20'h0bb4a: out <= 12'h088;
      20'h0bb4b: out <= 12'h088;
      20'h0bb4c: out <= 12'h088;
      20'h0bb4d: out <= 12'h088;
      20'h0bb4e: out <= 12'h088;
      20'h0bb4f: out <= 12'h088;
      20'h0bb50: out <= 12'h088;
      20'h0bb51: out <= 12'h088;
      20'h0bb52: out <= 12'h088;
      20'h0bb53: out <= 12'h088;
      20'h0bb54: out <= 12'h088;
      20'h0bb55: out <= 12'h088;
      20'h0bb56: out <= 12'h088;
      20'h0bb57: out <= 12'h088;
      20'h0bb58: out <= 12'h088;
      20'h0bb59: out <= 12'h088;
      20'h0bb5a: out <= 12'h088;
      20'h0bb5b: out <= 12'h088;
      20'h0bb5c: out <= 12'h088;
      20'h0bb5d: out <= 12'h088;
      20'h0bb5e: out <= 12'h088;
      20'h0bb5f: out <= 12'h088;
      20'h0bb60: out <= 12'h088;
      20'h0bb61: out <= 12'h088;
      20'h0bb62: out <= 12'h088;
      20'h0bb63: out <= 12'h088;
      20'h0bb64: out <= 12'h088;
      20'h0bb65: out <= 12'h088;
      20'h0bb66: out <= 12'h088;
      20'h0bb67: out <= 12'h088;
      20'h0bb68: out <= 12'h088;
      20'h0bb69: out <= 12'h088;
      20'h0bb6a: out <= 12'h088;
      20'h0bb6b: out <= 12'h088;
      20'h0bb6c: out <= 12'h088;
      20'h0bb6d: out <= 12'h088;
      20'h0bb6e: out <= 12'h088;
      20'h0bb6f: out <= 12'h088;
      20'h0bb70: out <= 12'h088;
      20'h0bb71: out <= 12'h222;
      20'h0bb72: out <= 12'h222;
      20'h0bb73: out <= 12'h222;
      20'h0bb74: out <= 12'h222;
      20'h0bb75: out <= 12'h222;
      20'h0bb76: out <= 12'h222;
      20'h0bb77: out <= 12'h222;
      20'h0bb78: out <= 12'h660;
      20'h0bb79: out <= 12'hbb0;
      20'h0bb7a: out <= 12'hee9;
      20'h0bb7b: out <= 12'hee9;
      20'h0bb7c: out <= 12'hee9;
      20'h0bb7d: out <= 12'hee9;
      20'h0bb7e: out <= 12'hee9;
      20'h0bb7f: out <= 12'hbb0;
      20'h0bb80: out <= 12'h660;
      20'h0bb81: out <= 12'h222;
      20'h0bb82: out <= 12'h222;
      20'h0bb83: out <= 12'h222;
      20'h0bb84: out <= 12'h222;
      20'h0bb85: out <= 12'h222;
      20'h0bb86: out <= 12'h222;
      20'h0bb87: out <= 12'h222;
      20'h0bb88: out <= 12'h603;
      20'h0bb89: out <= 12'h603;
      20'h0bb8a: out <= 12'h603;
      20'h0bb8b: out <= 12'h603;
      20'h0bb8c: out <= 12'hf87;
      20'h0bb8d: out <= 12'hf87;
      20'h0bb8e: out <= 12'h000;
      20'h0bb8f: out <= 12'h000;
      20'h0bb90: out <= 12'h000;
      20'h0bb91: out <= 12'hf87;
      20'h0bb92: out <= 12'hf87;
      20'h0bb93: out <= 12'h000;
      20'h0bb94: out <= 12'h000;
      20'h0bb95: out <= 12'h000;
      20'h0bb96: out <= 12'hf87;
      20'h0bb97: out <= 12'hf87;
      20'h0bb98: out <= 12'hf87;
      20'h0bb99: out <= 12'h000;
      20'h0bb9a: out <= 12'h000;
      20'h0bb9b: out <= 12'h000;
      20'h0bb9c: out <= 12'hf87;
      20'h0bb9d: out <= 12'hf87;
      20'h0bb9e: out <= 12'h000;
      20'h0bb9f: out <= 12'h000;
      20'h0bba0: out <= 12'h000;
      20'h0bba1: out <= 12'hf87;
      20'h0bba2: out <= 12'hf87;
      20'h0bba3: out <= 12'h000;
      20'h0bba4: out <= 12'hf87;
      20'h0bba5: out <= 12'hf87;
      20'h0bba6: out <= 12'h000;
      20'h0bba7: out <= 12'h000;
      20'h0bba8: out <= 12'h000;
      20'h0bba9: out <= 12'hf87;
      20'h0bbaa: out <= 12'hf87;
      20'h0bbab: out <= 12'h000;
      20'h0bbac: out <= 12'h000;
      20'h0bbad: out <= 12'h000;
      20'h0bbae: out <= 12'hf87;
      20'h0bbaf: out <= 12'hf87;
      20'h0bbb0: out <= 12'hf87;
      20'h0bbb1: out <= 12'hf87;
      20'h0bbb2: out <= 12'h000;
      20'h0bbb3: out <= 12'h000;
      20'h0bbb4: out <= 12'hf87;
      20'h0bbb5: out <= 12'hf87;
      20'h0bbb6: out <= 12'h000;
      20'h0bbb7: out <= 12'h000;
      20'h0bbb8: out <= 12'h000;
      20'h0bbb9: out <= 12'h000;
      20'h0bbba: out <= 12'h000;
      20'h0bbbb: out <= 12'h000;
      20'h0bbbc: out <= 12'hf87;
      20'h0bbbd: out <= 12'hf87;
      20'h0bbbe: out <= 12'hf87;
      20'h0bbbf: out <= 12'h000;
      20'h0bbc0: out <= 12'h000;
      20'h0bbc1: out <= 12'h000;
      20'h0bbc2: out <= 12'h000;
      20'h0bbc3: out <= 12'h000;
      20'h0bbc4: out <= 12'hf87;
      20'h0bbc5: out <= 12'hf87;
      20'h0bbc6: out <= 12'h000;
      20'h0bbc7: out <= 12'h000;
      20'h0bbc8: out <= 12'h000;
      20'h0bbc9: out <= 12'hf87;
      20'h0bbca: out <= 12'hf87;
      20'h0bbcb: out <= 12'h000;
      20'h0bbcc: out <= 12'hf87;
      20'h0bbcd: out <= 12'hf87;
      20'h0bbce: out <= 12'h000;
      20'h0bbcf: out <= 12'h000;
      20'h0bbd0: out <= 12'h000;
      20'h0bbd1: out <= 12'hf87;
      20'h0bbd2: out <= 12'hf87;
      20'h0bbd3: out <= 12'h000;
      20'h0bbd4: out <= 12'hf87;
      20'h0bbd5: out <= 12'hf87;
      20'h0bbd6: out <= 12'h000;
      20'h0bbd7: out <= 12'h000;
      20'h0bbd8: out <= 12'h000;
      20'h0bbd9: out <= 12'hf87;
      20'h0bbda: out <= 12'hf87;
      20'h0bbdb: out <= 12'h000;
      20'h0bbdc: out <= 12'h603;
      20'h0bbdd: out <= 12'h603;
      20'h0bbde: out <= 12'h603;
      20'h0bbdf: out <= 12'h603;
      20'h0bbe0: out <= 12'hee9;
      20'h0bbe1: out <= 12'hf87;
      20'h0bbe2: out <= 12'hee9;
      20'h0bbe3: out <= 12'hf87;
      20'h0bbe4: out <= 12'hf87;
      20'h0bbe5: out <= 12'hb27;
      20'h0bbe6: out <= 12'hf87;
      20'h0bbe7: out <= 12'hb27;
      20'h0bbe8: out <= 12'h000;
      20'h0bbe9: out <= 12'h000;
      20'h0bbea: out <= 12'h000;
      20'h0bbeb: out <= 12'h000;
      20'h0bbec: out <= 12'h000;
      20'h0bbed: out <= 12'h000;
      20'h0bbee: out <= 12'h000;
      20'h0bbef: out <= 12'h000;
      20'h0bbf0: out <= 12'h777;
      20'h0bbf1: out <= 12'h555;
      20'h0bbf2: out <= 12'h555;
      20'h0bbf3: out <= 12'h555;
      20'h0bbf4: out <= 12'h555;
      20'h0bbf5: out <= 12'h555;
      20'h0bbf6: out <= 12'h555;
      20'h0bbf7: out <= 12'h555;
      20'h0bbf8: out <= 12'h555;
      20'h0bbf9: out <= 12'h555;
      20'h0bbfa: out <= 12'h555;
      20'h0bbfb: out <= 12'h555;
      20'h0bbfc: out <= 12'h555;
      20'h0bbfd: out <= 12'h555;
      20'h0bbfe: out <= 12'h555;
      20'h0bbff: out <= 12'h777;
      20'h0bc00: out <= 12'h000;
      20'h0bc01: out <= 12'h000;
      20'h0bc02: out <= 12'h000;
      20'h0bc03: out <= 12'h000;
      20'h0bc04: out <= 12'hf87;
      20'h0bc05: out <= 12'h000;
      20'h0bc06: out <= 12'h000;
      20'h0bc07: out <= 12'h000;
      20'h0bc08: out <= 12'hfa9;
      20'h0bc09: out <= 12'hfa9;
      20'h0bc0a: out <= 12'hfa9;
      20'h0bc0b: out <= 12'hfa9;
      20'h0bc0c: out <= 12'hfa9;
      20'h0bc0d: out <= 12'hfa9;
      20'h0bc0e: out <= 12'hfa9;
      20'h0bc0f: out <= 12'hfa9;
      20'h0bc10: out <= 12'hf76;
      20'h0bc11: out <= 12'hf76;
      20'h0bc12: out <= 12'hf76;
      20'h0bc13: out <= 12'hf76;
      20'h0bc14: out <= 12'hf76;
      20'h0bc15: out <= 12'hf76;
      20'h0bc16: out <= 12'hf76;
      20'h0bc17: out <= 12'hf76;
      20'h0bc18: out <= 12'h000;
      20'h0bc19: out <= 12'h000;
      20'h0bc1a: out <= 12'h000;
      20'h0bc1b: out <= 12'h000;
      20'h0bc1c: out <= 12'h000;
      20'h0bc1d: out <= 12'h000;
      20'h0bc1e: out <= 12'h000;
      20'h0bc1f: out <= 12'h000;
      20'h0bc20: out <= 12'h088;
      20'h0bc21: out <= 12'h088;
      20'h0bc22: out <= 12'h088;
      20'h0bc23: out <= 12'h088;
      20'h0bc24: out <= 12'h088;
      20'h0bc25: out <= 12'h088;
      20'h0bc26: out <= 12'h088;
      20'h0bc27: out <= 12'h088;
      20'h0bc28: out <= 12'h088;
      20'h0bc29: out <= 12'h088;
      20'h0bc2a: out <= 12'h088;
      20'h0bc2b: out <= 12'h088;
      20'h0bc2c: out <= 12'h088;
      20'h0bc2d: out <= 12'h088;
      20'h0bc2e: out <= 12'h088;
      20'h0bc2f: out <= 12'h088;
      20'h0bc30: out <= 12'h088;
      20'h0bc31: out <= 12'h088;
      20'h0bc32: out <= 12'h088;
      20'h0bc33: out <= 12'h088;
      20'h0bc34: out <= 12'h088;
      20'h0bc35: out <= 12'h088;
      20'h0bc36: out <= 12'h088;
      20'h0bc37: out <= 12'h088;
      20'h0bc38: out <= 12'h088;
      20'h0bc39: out <= 12'h088;
      20'h0bc3a: out <= 12'h088;
      20'h0bc3b: out <= 12'h088;
      20'h0bc3c: out <= 12'h088;
      20'h0bc3d: out <= 12'h088;
      20'h0bc3e: out <= 12'h088;
      20'h0bc3f: out <= 12'h088;
      20'h0bc40: out <= 12'h088;
      20'h0bc41: out <= 12'h088;
      20'h0bc42: out <= 12'h088;
      20'h0bc43: out <= 12'h088;
      20'h0bc44: out <= 12'h088;
      20'h0bc45: out <= 12'h088;
      20'h0bc46: out <= 12'h088;
      20'h0bc47: out <= 12'h088;
      20'h0bc48: out <= 12'h088;
      20'h0bc49: out <= 12'h088;
      20'h0bc4a: out <= 12'h088;
      20'h0bc4b: out <= 12'h088;
      20'h0bc4c: out <= 12'h088;
      20'h0bc4d: out <= 12'h088;
      20'h0bc4e: out <= 12'h088;
      20'h0bc4f: out <= 12'h088;
      20'h0bc50: out <= 12'h088;
      20'h0bc51: out <= 12'h088;
      20'h0bc52: out <= 12'h088;
      20'h0bc53: out <= 12'h088;
      20'h0bc54: out <= 12'h088;
      20'h0bc55: out <= 12'h088;
      20'h0bc56: out <= 12'h088;
      20'h0bc57: out <= 12'h088;
      20'h0bc58: out <= 12'h088;
      20'h0bc59: out <= 12'h088;
      20'h0bc5a: out <= 12'h088;
      20'h0bc5b: out <= 12'h088;
      20'h0bc5c: out <= 12'h088;
      20'h0bc5d: out <= 12'h088;
      20'h0bc5e: out <= 12'h088;
      20'h0bc5f: out <= 12'h088;
      20'h0bc60: out <= 12'h088;
      20'h0bc61: out <= 12'h088;
      20'h0bc62: out <= 12'h088;
      20'h0bc63: out <= 12'h088;
      20'h0bc64: out <= 12'h088;
      20'h0bc65: out <= 12'h088;
      20'h0bc66: out <= 12'h088;
      20'h0bc67: out <= 12'h088;
      20'h0bc68: out <= 12'h088;
      20'h0bc69: out <= 12'h088;
      20'h0bc6a: out <= 12'h088;
      20'h0bc6b: out <= 12'h088;
      20'h0bc6c: out <= 12'h088;
      20'h0bc6d: out <= 12'h088;
      20'h0bc6e: out <= 12'h088;
      20'h0bc6f: out <= 12'h088;
      20'h0bc70: out <= 12'h088;
      20'h0bc71: out <= 12'h088;
      20'h0bc72: out <= 12'h088;
      20'h0bc73: out <= 12'h088;
      20'h0bc74: out <= 12'h088;
      20'h0bc75: out <= 12'h088;
      20'h0bc76: out <= 12'h088;
      20'h0bc77: out <= 12'h088;
      20'h0bc78: out <= 12'h088;
      20'h0bc79: out <= 12'h088;
      20'h0bc7a: out <= 12'h088;
      20'h0bc7b: out <= 12'h088;
      20'h0bc7c: out <= 12'h088;
      20'h0bc7d: out <= 12'h088;
      20'h0bc7e: out <= 12'h088;
      20'h0bc7f: out <= 12'h088;
      20'h0bc80: out <= 12'h088;
      20'h0bc81: out <= 12'h088;
      20'h0bc82: out <= 12'h088;
      20'h0bc83: out <= 12'h088;
      20'h0bc84: out <= 12'h088;
      20'h0bc85: out <= 12'h088;
      20'h0bc86: out <= 12'h088;
      20'h0bc87: out <= 12'h088;
      20'h0bc88: out <= 12'h088;
      20'h0bc89: out <= 12'h222;
      20'h0bc8a: out <= 12'h222;
      20'h0bc8b: out <= 12'h222;
      20'h0bc8c: out <= 12'h222;
      20'h0bc8d: out <= 12'h222;
      20'h0bc8e: out <= 12'h222;
      20'h0bc8f: out <= 12'h660;
      20'h0bc90: out <= 12'hbb0;
      20'h0bc91: out <= 12'hee9;
      20'h0bc92: out <= 12'hee9;
      20'h0bc93: out <= 12'hee9;
      20'h0bc94: out <= 12'hee9;
      20'h0bc95: out <= 12'hee9;
      20'h0bc96: out <= 12'hee9;
      20'h0bc97: out <= 12'hee9;
      20'h0bc98: out <= 12'hbb0;
      20'h0bc99: out <= 12'h660;
      20'h0bc9a: out <= 12'h222;
      20'h0bc9b: out <= 12'h222;
      20'h0bc9c: out <= 12'h222;
      20'h0bc9d: out <= 12'h222;
      20'h0bc9e: out <= 12'h222;
      20'h0bc9f: out <= 12'h222;
      20'h0bca0: out <= 12'h603;
      20'h0bca1: out <= 12'h603;
      20'h0bca2: out <= 12'h603;
      20'h0bca3: out <= 12'h603;
      20'h0bca4: out <= 12'hee9;
      20'h0bca5: out <= 12'hee9;
      20'h0bca6: out <= 12'h000;
      20'h0bca7: out <= 12'h000;
      20'h0bca8: out <= 12'hee9;
      20'h0bca9: out <= 12'hee9;
      20'h0bcaa: out <= 12'hee9;
      20'h0bcab: out <= 12'h000;
      20'h0bcac: out <= 12'h000;
      20'h0bcad: out <= 12'h000;
      20'h0bcae: out <= 12'h000;
      20'h0bcaf: out <= 12'hee9;
      20'h0bcb0: out <= 12'hee9;
      20'h0bcb1: out <= 12'h000;
      20'h0bcb2: out <= 12'h000;
      20'h0bcb3: out <= 12'h000;
      20'h0bcb4: out <= 12'h000;
      20'h0bcb5: out <= 12'h000;
      20'h0bcb6: out <= 12'h000;
      20'h0bcb7: out <= 12'h000;
      20'h0bcb8: out <= 12'h000;
      20'h0bcb9: out <= 12'hee9;
      20'h0bcba: out <= 12'hee9;
      20'h0bcbb: out <= 12'h000;
      20'h0bcbc: out <= 12'h000;
      20'h0bcbd: out <= 12'h000;
      20'h0bcbe: out <= 12'h000;
      20'h0bcbf: out <= 12'h000;
      20'h0bcc0: out <= 12'h000;
      20'h0bcc1: out <= 12'hee9;
      20'h0bcc2: out <= 12'hee9;
      20'h0bcc3: out <= 12'h000;
      20'h0bcc4: out <= 12'h000;
      20'h0bcc5: out <= 12'hee9;
      20'h0bcc6: out <= 12'hee9;
      20'h0bcc7: out <= 12'h000;
      20'h0bcc8: out <= 12'hee9;
      20'h0bcc9: out <= 12'hee9;
      20'h0bcca: out <= 12'h000;
      20'h0bccb: out <= 12'h000;
      20'h0bccc: out <= 12'hee9;
      20'h0bccd: out <= 12'hee9;
      20'h0bcce: out <= 12'h000;
      20'h0bccf: out <= 12'h000;
      20'h0bcd0: out <= 12'h000;
      20'h0bcd1: out <= 12'h000;
      20'h0bcd2: out <= 12'h000;
      20'h0bcd3: out <= 12'h000;
      20'h0bcd4: out <= 12'hee9;
      20'h0bcd5: out <= 12'hee9;
      20'h0bcd6: out <= 12'h000;
      20'h0bcd7: out <= 12'h000;
      20'h0bcd8: out <= 12'h000;
      20'h0bcd9: out <= 12'h000;
      20'h0bcda: out <= 12'h000;
      20'h0bcdb: out <= 12'h000;
      20'h0bcdc: out <= 12'h000;
      20'h0bcdd: out <= 12'h000;
      20'h0bcde: out <= 12'h000;
      20'h0bcdf: out <= 12'h000;
      20'h0bce0: out <= 12'h000;
      20'h0bce1: out <= 12'hee9;
      20'h0bce2: out <= 12'hee9;
      20'h0bce3: out <= 12'h000;
      20'h0bce4: out <= 12'hee9;
      20'h0bce5: out <= 12'hee9;
      20'h0bce6: out <= 12'h000;
      20'h0bce7: out <= 12'h000;
      20'h0bce8: out <= 12'h000;
      20'h0bce9: out <= 12'hee9;
      20'h0bcea: out <= 12'hee9;
      20'h0bceb: out <= 12'h000;
      20'h0bcec: out <= 12'hee9;
      20'h0bced: out <= 12'hee9;
      20'h0bcee: out <= 12'h000;
      20'h0bcef: out <= 12'h000;
      20'h0bcf0: out <= 12'h000;
      20'h0bcf1: out <= 12'hee9;
      20'h0bcf2: out <= 12'hee9;
      20'h0bcf3: out <= 12'h000;
      20'h0bcf4: out <= 12'h603;
      20'h0bcf5: out <= 12'h603;
      20'h0bcf6: out <= 12'h603;
      20'h0bcf7: out <= 12'h603;
      20'h0bcf8: out <= 12'hee9;
      20'h0bcf9: out <= 12'hf87;
      20'h0bcfa: out <= 12'hee9;
      20'h0bcfb: out <= 12'hf87;
      20'h0bcfc: out <= 12'hf87;
      20'h0bcfd: out <= 12'hb27;
      20'h0bcfe: out <= 12'hf87;
      20'h0bcff: out <= 12'hb27;
      20'h0bd00: out <= 12'h000;
      20'h0bd01: out <= 12'h000;
      20'h0bd02: out <= 12'h000;
      20'h0bd03: out <= 12'h000;
      20'h0bd04: out <= 12'h000;
      20'h0bd05: out <= 12'h000;
      20'h0bd06: out <= 12'h000;
      20'h0bd07: out <= 12'h000;
      20'h0bd08: out <= 12'h777;
      20'h0bd09: out <= 12'h555;
      20'h0bd0a: out <= 12'h555;
      20'h0bd0b: out <= 12'h555;
      20'h0bd0c: out <= 12'h555;
      20'h0bd0d: out <= 12'h555;
      20'h0bd0e: out <= 12'h555;
      20'h0bd0f: out <= 12'h555;
      20'h0bd10: out <= 12'h555;
      20'h0bd11: out <= 12'h555;
      20'h0bd12: out <= 12'h555;
      20'h0bd13: out <= 12'h555;
      20'h0bd14: out <= 12'h555;
      20'h0bd15: out <= 12'h555;
      20'h0bd16: out <= 12'h555;
      20'h0bd17: out <= 12'h777;
      20'h0bd18: out <= 12'h000;
      20'h0bd19: out <= 12'h000;
      20'h0bd1a: out <= 12'h000;
      20'h0bd1b: out <= 12'hf87;
      20'h0bd1c: out <= 12'h000;
      20'h0bd1d: out <= 12'hf87;
      20'h0bd1e: out <= 12'h000;
      20'h0bd1f: out <= 12'h000;
      20'h0bd20: out <= 12'hfa9;
      20'h0bd21: out <= 12'hfa9;
      20'h0bd22: out <= 12'hfa9;
      20'h0bd23: out <= 12'hfa9;
      20'h0bd24: out <= 12'hfa9;
      20'h0bd25: out <= 12'hfa9;
      20'h0bd26: out <= 12'hfa9;
      20'h0bd27: out <= 12'hfa9;
      20'h0bd28: out <= 12'hf76;
      20'h0bd29: out <= 12'hf76;
      20'h0bd2a: out <= 12'hf76;
      20'h0bd2b: out <= 12'hf76;
      20'h0bd2c: out <= 12'hf76;
      20'h0bd2d: out <= 12'hf76;
      20'h0bd2e: out <= 12'hf76;
      20'h0bd2f: out <= 12'hf76;
      20'h0bd30: out <= 12'h000;
      20'h0bd31: out <= 12'h000;
      20'h0bd32: out <= 12'h000;
      20'h0bd33: out <= 12'h000;
      20'h0bd34: out <= 12'h000;
      20'h0bd35: out <= 12'h000;
      20'h0bd36: out <= 12'h000;
      20'h0bd37: out <= 12'h000;
      20'h0bd38: out <= 12'h088;
      20'h0bd39: out <= 12'h088;
      20'h0bd3a: out <= 12'h088;
      20'h0bd3b: out <= 12'h088;
      20'h0bd3c: out <= 12'h088;
      20'h0bd3d: out <= 12'h088;
      20'h0bd3e: out <= 12'h088;
      20'h0bd3f: out <= 12'h088;
      20'h0bd40: out <= 12'h088;
      20'h0bd41: out <= 12'h088;
      20'h0bd42: out <= 12'h088;
      20'h0bd43: out <= 12'h088;
      20'h0bd44: out <= 12'h088;
      20'h0bd45: out <= 12'h088;
      20'h0bd46: out <= 12'h088;
      20'h0bd47: out <= 12'h088;
      20'h0bd48: out <= 12'h088;
      20'h0bd49: out <= 12'h088;
      20'h0bd4a: out <= 12'h088;
      20'h0bd4b: out <= 12'h088;
      20'h0bd4c: out <= 12'h088;
      20'h0bd4d: out <= 12'h088;
      20'h0bd4e: out <= 12'h088;
      20'h0bd4f: out <= 12'h088;
      20'h0bd50: out <= 12'h088;
      20'h0bd51: out <= 12'h088;
      20'h0bd52: out <= 12'h088;
      20'h0bd53: out <= 12'h088;
      20'h0bd54: out <= 12'h088;
      20'h0bd55: out <= 12'h088;
      20'h0bd56: out <= 12'h088;
      20'h0bd57: out <= 12'h088;
      20'h0bd58: out <= 12'h088;
      20'h0bd59: out <= 12'h088;
      20'h0bd5a: out <= 12'h088;
      20'h0bd5b: out <= 12'h088;
      20'h0bd5c: out <= 12'h088;
      20'h0bd5d: out <= 12'h088;
      20'h0bd5e: out <= 12'h088;
      20'h0bd5f: out <= 12'h088;
      20'h0bd60: out <= 12'h088;
      20'h0bd61: out <= 12'h088;
      20'h0bd62: out <= 12'h088;
      20'h0bd63: out <= 12'h088;
      20'h0bd64: out <= 12'h088;
      20'h0bd65: out <= 12'h088;
      20'h0bd66: out <= 12'h088;
      20'h0bd67: out <= 12'h088;
      20'h0bd68: out <= 12'h088;
      20'h0bd69: out <= 12'h088;
      20'h0bd6a: out <= 12'h088;
      20'h0bd6b: out <= 12'h088;
      20'h0bd6c: out <= 12'h088;
      20'h0bd6d: out <= 12'h088;
      20'h0bd6e: out <= 12'h088;
      20'h0bd6f: out <= 12'h088;
      20'h0bd70: out <= 12'h088;
      20'h0bd71: out <= 12'h088;
      20'h0bd72: out <= 12'h088;
      20'h0bd73: out <= 12'h088;
      20'h0bd74: out <= 12'h088;
      20'h0bd75: out <= 12'h088;
      20'h0bd76: out <= 12'h088;
      20'h0bd77: out <= 12'h088;
      20'h0bd78: out <= 12'h088;
      20'h0bd79: out <= 12'h088;
      20'h0bd7a: out <= 12'h088;
      20'h0bd7b: out <= 12'h088;
      20'h0bd7c: out <= 12'h088;
      20'h0bd7d: out <= 12'h088;
      20'h0bd7e: out <= 12'h088;
      20'h0bd7f: out <= 12'h088;
      20'h0bd80: out <= 12'h088;
      20'h0bd81: out <= 12'h088;
      20'h0bd82: out <= 12'h088;
      20'h0bd83: out <= 12'h088;
      20'h0bd84: out <= 12'h088;
      20'h0bd85: out <= 12'h088;
      20'h0bd86: out <= 12'h088;
      20'h0bd87: out <= 12'h088;
      20'h0bd88: out <= 12'h088;
      20'h0bd89: out <= 12'h088;
      20'h0bd8a: out <= 12'h088;
      20'h0bd8b: out <= 12'h088;
      20'h0bd8c: out <= 12'h088;
      20'h0bd8d: out <= 12'h088;
      20'h0bd8e: out <= 12'h088;
      20'h0bd8f: out <= 12'h088;
      20'h0bd90: out <= 12'h088;
      20'h0bd91: out <= 12'h088;
      20'h0bd92: out <= 12'h088;
      20'h0bd93: out <= 12'h088;
      20'h0bd94: out <= 12'h088;
      20'h0bd95: out <= 12'h088;
      20'h0bd96: out <= 12'h088;
      20'h0bd97: out <= 12'h088;
      20'h0bd98: out <= 12'h088;
      20'h0bd99: out <= 12'h088;
      20'h0bd9a: out <= 12'h088;
      20'h0bd9b: out <= 12'h088;
      20'h0bd9c: out <= 12'h088;
      20'h0bd9d: out <= 12'h088;
      20'h0bd9e: out <= 12'h088;
      20'h0bd9f: out <= 12'h088;
      20'h0bda0: out <= 12'h088;
      20'h0bda1: out <= 12'h222;
      20'h0bda2: out <= 12'h222;
      20'h0bda3: out <= 12'h222;
      20'h0bda4: out <= 12'h222;
      20'h0bda5: out <= 12'h222;
      20'h0bda6: out <= 12'h660;
      20'h0bda7: out <= 12'hbb0;
      20'h0bda8: out <= 12'hee9;
      20'h0bda9: out <= 12'hee9;
      20'h0bdaa: out <= 12'hee9;
      20'h0bdab: out <= 12'hee9;
      20'h0bdac: out <= 12'hee9;
      20'h0bdad: out <= 12'hee9;
      20'h0bdae: out <= 12'hee9;
      20'h0bdaf: out <= 12'hee9;
      20'h0bdb0: out <= 12'hee9;
      20'h0bdb1: out <= 12'hbb0;
      20'h0bdb2: out <= 12'h660;
      20'h0bdb3: out <= 12'h222;
      20'h0bdb4: out <= 12'h222;
      20'h0bdb5: out <= 12'h222;
      20'h0bdb6: out <= 12'h222;
      20'h0bdb7: out <= 12'h222;
      20'h0bdb8: out <= 12'h603;
      20'h0bdb9: out <= 12'h603;
      20'h0bdba: out <= 12'h603;
      20'h0bdbb: out <= 12'h603;
      20'h0bdbc: out <= 12'hee9;
      20'h0bdbd: out <= 12'hee9;
      20'h0bdbe: out <= 12'h000;
      20'h0bdbf: out <= 12'h000;
      20'h0bdc0: out <= 12'hee9;
      20'h0bdc1: out <= 12'hee9;
      20'h0bdc2: out <= 12'hee9;
      20'h0bdc3: out <= 12'h000;
      20'h0bdc4: out <= 12'h000;
      20'h0bdc5: out <= 12'h000;
      20'h0bdc6: out <= 12'h000;
      20'h0bdc7: out <= 12'hee9;
      20'h0bdc8: out <= 12'hee9;
      20'h0bdc9: out <= 12'h000;
      20'h0bdca: out <= 12'h000;
      20'h0bdcb: out <= 12'h000;
      20'h0bdcc: out <= 12'h000;
      20'h0bdcd: out <= 12'h000;
      20'h0bdce: out <= 12'h000;
      20'h0bdcf: out <= 12'h000;
      20'h0bdd0: out <= 12'hee9;
      20'h0bdd1: out <= 12'hee9;
      20'h0bdd2: out <= 12'hee9;
      20'h0bdd3: out <= 12'h000;
      20'h0bdd4: out <= 12'h000;
      20'h0bdd5: out <= 12'h000;
      20'h0bdd6: out <= 12'h000;
      20'h0bdd7: out <= 12'h000;
      20'h0bdd8: out <= 12'h000;
      20'h0bdd9: out <= 12'hee9;
      20'h0bdda: out <= 12'hee9;
      20'h0bddb: out <= 12'h000;
      20'h0bddc: out <= 12'h000;
      20'h0bddd: out <= 12'hee9;
      20'h0bdde: out <= 12'hee9;
      20'h0bddf: out <= 12'h000;
      20'h0bde0: out <= 12'hee9;
      20'h0bde1: out <= 12'hee9;
      20'h0bde2: out <= 12'h000;
      20'h0bde3: out <= 12'h000;
      20'h0bde4: out <= 12'hee9;
      20'h0bde5: out <= 12'hee9;
      20'h0bde6: out <= 12'hee9;
      20'h0bde7: out <= 12'hee9;
      20'h0bde8: out <= 12'hee9;
      20'h0bde9: out <= 12'hee9;
      20'h0bdea: out <= 12'h000;
      20'h0bdeb: out <= 12'h000;
      20'h0bdec: out <= 12'hee9;
      20'h0bded: out <= 12'hee9;
      20'h0bdee: out <= 12'h000;
      20'h0bdef: out <= 12'h000;
      20'h0bdf0: out <= 12'h000;
      20'h0bdf1: out <= 12'h000;
      20'h0bdf2: out <= 12'h000;
      20'h0bdf3: out <= 12'h000;
      20'h0bdf4: out <= 12'h000;
      20'h0bdf5: out <= 12'h000;
      20'h0bdf6: out <= 12'h000;
      20'h0bdf7: out <= 12'h000;
      20'h0bdf8: out <= 12'hee9;
      20'h0bdf9: out <= 12'hee9;
      20'h0bdfa: out <= 12'h000;
      20'h0bdfb: out <= 12'h000;
      20'h0bdfc: out <= 12'hee9;
      20'h0bdfd: out <= 12'hee9;
      20'h0bdfe: out <= 12'h000;
      20'h0bdff: out <= 12'h000;
      20'h0be00: out <= 12'h000;
      20'h0be01: out <= 12'hee9;
      20'h0be02: out <= 12'hee9;
      20'h0be03: out <= 12'h000;
      20'h0be04: out <= 12'hee9;
      20'h0be05: out <= 12'hee9;
      20'h0be06: out <= 12'h000;
      20'h0be07: out <= 12'h000;
      20'h0be08: out <= 12'h000;
      20'h0be09: out <= 12'hee9;
      20'h0be0a: out <= 12'hee9;
      20'h0be0b: out <= 12'h000;
      20'h0be0c: out <= 12'h603;
      20'h0be0d: out <= 12'h603;
      20'h0be0e: out <= 12'h603;
      20'h0be0f: out <= 12'h603;
      20'h0be10: out <= 12'hee9;
      20'h0be11: out <= 12'hf87;
      20'h0be12: out <= 12'hee9;
      20'h0be13: out <= 12'hb27;
      20'h0be14: out <= 12'hb27;
      20'h0be15: out <= 12'hb27;
      20'h0be16: out <= 12'hf87;
      20'h0be17: out <= 12'hb27;
      20'h0be18: out <= 12'h000;
      20'h0be19: out <= 12'h000;
      20'h0be1a: out <= 12'h000;
      20'h0be1b: out <= 12'h000;
      20'h0be1c: out <= 12'h000;
      20'h0be1d: out <= 12'h000;
      20'h0be1e: out <= 12'h000;
      20'h0be1f: out <= 12'h000;
      20'h0be20: out <= 12'h777;
      20'h0be21: out <= 12'h555;
      20'h0be22: out <= 12'h555;
      20'h0be23: out <= 12'h555;
      20'h0be24: out <= 12'h555;
      20'h0be25: out <= 12'h555;
      20'h0be26: out <= 12'h555;
      20'h0be27: out <= 12'h555;
      20'h0be28: out <= 12'h555;
      20'h0be29: out <= 12'h555;
      20'h0be2a: out <= 12'h555;
      20'h0be2b: out <= 12'h555;
      20'h0be2c: out <= 12'h555;
      20'h0be2d: out <= 12'h555;
      20'h0be2e: out <= 12'h555;
      20'h0be2f: out <= 12'h777;
      20'h0be30: out <= 12'h000;
      20'h0be31: out <= 12'h000;
      20'h0be32: out <= 12'hf87;
      20'h0be33: out <= 12'h000;
      20'h0be34: out <= 12'h000;
      20'h0be35: out <= 12'h000;
      20'h0be36: out <= 12'hf87;
      20'h0be37: out <= 12'h000;
      20'h0be38: out <= 12'hfa9;
      20'h0be39: out <= 12'hfa9;
      20'h0be3a: out <= 12'hfa9;
      20'h0be3b: out <= 12'hfa9;
      20'h0be3c: out <= 12'hfa9;
      20'h0be3d: out <= 12'hfa9;
      20'h0be3e: out <= 12'hfa9;
      20'h0be3f: out <= 12'hfa9;
      20'h0be40: out <= 12'hf76;
      20'h0be41: out <= 12'hf76;
      20'h0be42: out <= 12'hf76;
      20'h0be43: out <= 12'hf76;
      20'h0be44: out <= 12'hf76;
      20'h0be45: out <= 12'hf76;
      20'h0be46: out <= 12'hf76;
      20'h0be47: out <= 12'hf76;
      20'h0be48: out <= 12'h000;
      20'h0be49: out <= 12'h000;
      20'h0be4a: out <= 12'h000;
      20'h0be4b: out <= 12'h000;
      20'h0be4c: out <= 12'h000;
      20'h0be4d: out <= 12'h000;
      20'h0be4e: out <= 12'h000;
      20'h0be4f: out <= 12'h000;
      20'h0be50: out <= 12'h088;
      20'h0be51: out <= 12'h088;
      20'h0be52: out <= 12'h088;
      20'h0be53: out <= 12'h088;
      20'h0be54: out <= 12'h088;
      20'h0be55: out <= 12'h088;
      20'h0be56: out <= 12'h088;
      20'h0be57: out <= 12'h088;
      20'h0be58: out <= 12'h088;
      20'h0be59: out <= 12'h088;
      20'h0be5a: out <= 12'h088;
      20'h0be5b: out <= 12'h088;
      20'h0be5c: out <= 12'h088;
      20'h0be5d: out <= 12'h088;
      20'h0be5e: out <= 12'h088;
      20'h0be5f: out <= 12'h088;
      20'h0be60: out <= 12'h088;
      20'h0be61: out <= 12'h088;
      20'h0be62: out <= 12'h088;
      20'h0be63: out <= 12'h088;
      20'h0be64: out <= 12'h088;
      20'h0be65: out <= 12'h088;
      20'h0be66: out <= 12'h088;
      20'h0be67: out <= 12'h088;
      20'h0be68: out <= 12'h088;
      20'h0be69: out <= 12'h088;
      20'h0be6a: out <= 12'h088;
      20'h0be6b: out <= 12'h088;
      20'h0be6c: out <= 12'h088;
      20'h0be6d: out <= 12'h088;
      20'h0be6e: out <= 12'h088;
      20'h0be6f: out <= 12'h088;
      20'h0be70: out <= 12'h088;
      20'h0be71: out <= 12'h088;
      20'h0be72: out <= 12'h088;
      20'h0be73: out <= 12'h088;
      20'h0be74: out <= 12'h088;
      20'h0be75: out <= 12'h088;
      20'h0be76: out <= 12'h088;
      20'h0be77: out <= 12'h088;
      20'h0be78: out <= 12'h088;
      20'h0be79: out <= 12'h088;
      20'h0be7a: out <= 12'h088;
      20'h0be7b: out <= 12'h088;
      20'h0be7c: out <= 12'h088;
      20'h0be7d: out <= 12'h088;
      20'h0be7e: out <= 12'h088;
      20'h0be7f: out <= 12'h088;
      20'h0be80: out <= 12'h088;
      20'h0be81: out <= 12'h088;
      20'h0be82: out <= 12'h088;
      20'h0be83: out <= 12'h088;
      20'h0be84: out <= 12'h088;
      20'h0be85: out <= 12'h088;
      20'h0be86: out <= 12'h088;
      20'h0be87: out <= 12'h088;
      20'h0be88: out <= 12'h088;
      20'h0be89: out <= 12'h088;
      20'h0be8a: out <= 12'h088;
      20'h0be8b: out <= 12'h088;
      20'h0be8c: out <= 12'h088;
      20'h0be8d: out <= 12'h088;
      20'h0be8e: out <= 12'h088;
      20'h0be8f: out <= 12'h088;
      20'h0be90: out <= 12'h088;
      20'h0be91: out <= 12'h088;
      20'h0be92: out <= 12'h088;
      20'h0be93: out <= 12'h088;
      20'h0be94: out <= 12'h088;
      20'h0be95: out <= 12'h088;
      20'h0be96: out <= 12'h088;
      20'h0be97: out <= 12'h088;
      20'h0be98: out <= 12'h088;
      20'h0be99: out <= 12'h088;
      20'h0be9a: out <= 12'h088;
      20'h0be9b: out <= 12'h088;
      20'h0be9c: out <= 12'h088;
      20'h0be9d: out <= 12'h088;
      20'h0be9e: out <= 12'h088;
      20'h0be9f: out <= 12'h088;
      20'h0bea0: out <= 12'h088;
      20'h0bea1: out <= 12'h088;
      20'h0bea2: out <= 12'h088;
      20'h0bea3: out <= 12'h088;
      20'h0bea4: out <= 12'h088;
      20'h0bea5: out <= 12'h088;
      20'h0bea6: out <= 12'h088;
      20'h0bea7: out <= 12'h088;
      20'h0bea8: out <= 12'h088;
      20'h0bea9: out <= 12'h088;
      20'h0beaa: out <= 12'h088;
      20'h0beab: out <= 12'h088;
      20'h0beac: out <= 12'h088;
      20'h0bead: out <= 12'h088;
      20'h0beae: out <= 12'h088;
      20'h0beaf: out <= 12'h088;
      20'h0beb0: out <= 12'h088;
      20'h0beb1: out <= 12'h088;
      20'h0beb2: out <= 12'h088;
      20'h0beb3: out <= 12'h088;
      20'h0beb4: out <= 12'h088;
      20'h0beb5: out <= 12'h088;
      20'h0beb6: out <= 12'h088;
      20'h0beb7: out <= 12'h088;
      20'h0beb8: out <= 12'h088;
      20'h0beb9: out <= 12'h222;
      20'h0beba: out <= 12'h222;
      20'h0bebb: out <= 12'h222;
      20'h0bebc: out <= 12'h222;
      20'h0bebd: out <= 12'h660;
      20'h0bebe: out <= 12'hbb0;
      20'h0bebf: out <= 12'hee9;
      20'h0bec0: out <= 12'hee9;
      20'h0bec1: out <= 12'hee9;
      20'h0bec2: out <= 12'hee9;
      20'h0bec3: out <= 12'hee9;
      20'h0bec4: out <= 12'hee9;
      20'h0bec5: out <= 12'hee9;
      20'h0bec6: out <= 12'hee9;
      20'h0bec7: out <= 12'hee9;
      20'h0bec8: out <= 12'hee9;
      20'h0bec9: out <= 12'hee9;
      20'h0beca: out <= 12'hbb0;
      20'h0becb: out <= 12'h660;
      20'h0becc: out <= 12'h222;
      20'h0becd: out <= 12'h222;
      20'h0bece: out <= 12'h222;
      20'h0becf: out <= 12'h222;
      20'h0bed0: out <= 12'h603;
      20'h0bed1: out <= 12'h603;
      20'h0bed2: out <= 12'h603;
      20'h0bed3: out <= 12'h603;
      20'h0bed4: out <= 12'hee9;
      20'h0bed5: out <= 12'hee9;
      20'h0bed6: out <= 12'h000;
      20'h0bed7: out <= 12'hee9;
      20'h0bed8: out <= 12'h000;
      20'h0bed9: out <= 12'hee9;
      20'h0beda: out <= 12'hee9;
      20'h0bedb: out <= 12'h000;
      20'h0bedc: out <= 12'h000;
      20'h0bedd: out <= 12'h000;
      20'h0bede: out <= 12'h000;
      20'h0bedf: out <= 12'hee9;
      20'h0bee0: out <= 12'hee9;
      20'h0bee1: out <= 12'h000;
      20'h0bee2: out <= 12'h000;
      20'h0bee3: out <= 12'h000;
      20'h0bee4: out <= 12'h000;
      20'h0bee5: out <= 12'h000;
      20'h0bee6: out <= 12'h000;
      20'h0bee7: out <= 12'h000;
      20'h0bee8: out <= 12'hee9;
      20'h0bee9: out <= 12'hee9;
      20'h0beea: out <= 12'h000;
      20'h0beeb: out <= 12'h000;
      20'h0beec: out <= 12'h000;
      20'h0beed: out <= 12'h000;
      20'h0beee: out <= 12'hee9;
      20'h0beef: out <= 12'hee9;
      20'h0bef0: out <= 12'hee9;
      20'h0bef1: out <= 12'hee9;
      20'h0bef2: out <= 12'h000;
      20'h0bef3: out <= 12'h000;
      20'h0bef4: out <= 12'h000;
      20'h0bef5: out <= 12'hee9;
      20'h0bef6: out <= 12'hee9;
      20'h0bef7: out <= 12'h000;
      20'h0bef8: out <= 12'hee9;
      20'h0bef9: out <= 12'hee9;
      20'h0befa: out <= 12'h000;
      20'h0befb: out <= 12'h000;
      20'h0befc: out <= 12'hee9;
      20'h0befd: out <= 12'hee9;
      20'h0befe: out <= 12'hee9;
      20'h0beff: out <= 12'hee9;
      20'h0bf00: out <= 12'hee9;
      20'h0bf01: out <= 12'hee9;
      20'h0bf02: out <= 12'hee9;
      20'h0bf03: out <= 12'h000;
      20'h0bf04: out <= 12'hee9;
      20'h0bf05: out <= 12'hee9;
      20'h0bf06: out <= 12'hee9;
      20'h0bf07: out <= 12'hee9;
      20'h0bf08: out <= 12'hee9;
      20'h0bf09: out <= 12'hee9;
      20'h0bf0a: out <= 12'h000;
      20'h0bf0b: out <= 12'h000;
      20'h0bf0c: out <= 12'h000;
      20'h0bf0d: out <= 12'h000;
      20'h0bf0e: out <= 12'h000;
      20'h0bf0f: out <= 12'h000;
      20'h0bf10: out <= 12'hee9;
      20'h0bf11: out <= 12'hee9;
      20'h0bf12: out <= 12'h000;
      20'h0bf13: out <= 12'h000;
      20'h0bf14: out <= 12'h000;
      20'h0bf15: out <= 12'hee9;
      20'h0bf16: out <= 12'hee9;
      20'h0bf17: out <= 12'hee9;
      20'h0bf18: out <= 12'hee9;
      20'h0bf19: out <= 12'hee9;
      20'h0bf1a: out <= 12'h000;
      20'h0bf1b: out <= 12'h000;
      20'h0bf1c: out <= 12'hee9;
      20'h0bf1d: out <= 12'hee9;
      20'h0bf1e: out <= 12'hee9;
      20'h0bf1f: out <= 12'hee9;
      20'h0bf20: out <= 12'hee9;
      20'h0bf21: out <= 12'hee9;
      20'h0bf22: out <= 12'hee9;
      20'h0bf23: out <= 12'h000;
      20'h0bf24: out <= 12'h603;
      20'h0bf25: out <= 12'h603;
      20'h0bf26: out <= 12'h603;
      20'h0bf27: out <= 12'h603;
      20'h0bf28: out <= 12'hee9;
      20'h0bf29: out <= 12'hf87;
      20'h0bf2a: out <= 12'hf87;
      20'h0bf2b: out <= 12'hf87;
      20'h0bf2c: out <= 12'hf87;
      20'h0bf2d: out <= 12'hf87;
      20'h0bf2e: out <= 12'hf87;
      20'h0bf2f: out <= 12'hb27;
      20'h0bf30: out <= 12'h000;
      20'h0bf31: out <= 12'h000;
      20'h0bf32: out <= 12'h000;
      20'h0bf33: out <= 12'h000;
      20'h0bf34: out <= 12'h000;
      20'h0bf35: out <= 12'h000;
      20'h0bf36: out <= 12'h000;
      20'h0bf37: out <= 12'h000;
      20'h0bf38: out <= 12'h777;
      20'h0bf39: out <= 12'h777;
      20'h0bf3a: out <= 12'h555;
      20'h0bf3b: out <= 12'h555;
      20'h0bf3c: out <= 12'h555;
      20'h0bf3d: out <= 12'h555;
      20'h0bf3e: out <= 12'h555;
      20'h0bf3f: out <= 12'h555;
      20'h0bf40: out <= 12'h555;
      20'h0bf41: out <= 12'h555;
      20'h0bf42: out <= 12'h555;
      20'h0bf43: out <= 12'h555;
      20'h0bf44: out <= 12'h555;
      20'h0bf45: out <= 12'h555;
      20'h0bf46: out <= 12'h777;
      20'h0bf47: out <= 12'h777;
      20'h0bf48: out <= 12'h000;
      20'h0bf49: out <= 12'h000;
      20'h0bf4a: out <= 12'h000;
      20'h0bf4b: out <= 12'h000;
      20'h0bf4c: out <= 12'h000;
      20'h0bf4d: out <= 12'h000;
      20'h0bf4e: out <= 12'h000;
      20'h0bf4f: out <= 12'h000;
      20'h0bf50: out <= 12'hfa9;
      20'h0bf51: out <= 12'hfa9;
      20'h0bf52: out <= 12'hfa9;
      20'h0bf53: out <= 12'hfa9;
      20'h0bf54: out <= 12'hfa9;
      20'h0bf55: out <= 12'hfa9;
      20'h0bf56: out <= 12'hfa9;
      20'h0bf57: out <= 12'hfa9;
      20'h0bf58: out <= 12'hf76;
      20'h0bf59: out <= 12'hf76;
      20'h0bf5a: out <= 12'hf76;
      20'h0bf5b: out <= 12'hf76;
      20'h0bf5c: out <= 12'hf76;
      20'h0bf5d: out <= 12'hf76;
      20'h0bf5e: out <= 12'hf76;
      20'h0bf5f: out <= 12'hf76;
      20'h0bf60: out <= 12'h000;
      20'h0bf61: out <= 12'h000;
      20'h0bf62: out <= 12'h000;
      20'h0bf63: out <= 12'h000;
      20'h0bf64: out <= 12'h000;
      20'h0bf65: out <= 12'h000;
      20'h0bf66: out <= 12'h000;
      20'h0bf67: out <= 12'h000;
      20'h0bf68: out <= 12'h088;
      20'h0bf69: out <= 12'h088;
      20'h0bf6a: out <= 12'h088;
      20'h0bf6b: out <= 12'h088;
      20'h0bf6c: out <= 12'h088;
      20'h0bf6d: out <= 12'h088;
      20'h0bf6e: out <= 12'h088;
      20'h0bf6f: out <= 12'h088;
      20'h0bf70: out <= 12'h088;
      20'h0bf71: out <= 12'h088;
      20'h0bf72: out <= 12'h088;
      20'h0bf73: out <= 12'h088;
      20'h0bf74: out <= 12'h088;
      20'h0bf75: out <= 12'h088;
      20'h0bf76: out <= 12'h088;
      20'h0bf77: out <= 12'h088;
      20'h0bf78: out <= 12'h088;
      20'h0bf79: out <= 12'h088;
      20'h0bf7a: out <= 12'h088;
      20'h0bf7b: out <= 12'h088;
      20'h0bf7c: out <= 12'h088;
      20'h0bf7d: out <= 12'h088;
      20'h0bf7e: out <= 12'h088;
      20'h0bf7f: out <= 12'h088;
      20'h0bf80: out <= 12'h088;
      20'h0bf81: out <= 12'h088;
      20'h0bf82: out <= 12'h088;
      20'h0bf83: out <= 12'h088;
      20'h0bf84: out <= 12'h088;
      20'h0bf85: out <= 12'h088;
      20'h0bf86: out <= 12'h088;
      20'h0bf87: out <= 12'h088;
      20'h0bf88: out <= 12'h088;
      20'h0bf89: out <= 12'h088;
      20'h0bf8a: out <= 12'h088;
      20'h0bf8b: out <= 12'h088;
      20'h0bf8c: out <= 12'h088;
      20'h0bf8d: out <= 12'h088;
      20'h0bf8e: out <= 12'h088;
      20'h0bf8f: out <= 12'h088;
      20'h0bf90: out <= 12'h088;
      20'h0bf91: out <= 12'h088;
      20'h0bf92: out <= 12'h088;
      20'h0bf93: out <= 12'h088;
      20'h0bf94: out <= 12'h088;
      20'h0bf95: out <= 12'h088;
      20'h0bf96: out <= 12'h088;
      20'h0bf97: out <= 12'h088;
      20'h0bf98: out <= 12'h088;
      20'h0bf99: out <= 12'h088;
      20'h0bf9a: out <= 12'h088;
      20'h0bf9b: out <= 12'h088;
      20'h0bf9c: out <= 12'h088;
      20'h0bf9d: out <= 12'h088;
      20'h0bf9e: out <= 12'h088;
      20'h0bf9f: out <= 12'h088;
      20'h0bfa0: out <= 12'h088;
      20'h0bfa1: out <= 12'h088;
      20'h0bfa2: out <= 12'h088;
      20'h0bfa3: out <= 12'h088;
      20'h0bfa4: out <= 12'h088;
      20'h0bfa5: out <= 12'h088;
      20'h0bfa6: out <= 12'h088;
      20'h0bfa7: out <= 12'h088;
      20'h0bfa8: out <= 12'h088;
      20'h0bfa9: out <= 12'h088;
      20'h0bfaa: out <= 12'h088;
      20'h0bfab: out <= 12'h088;
      20'h0bfac: out <= 12'h088;
      20'h0bfad: out <= 12'h088;
      20'h0bfae: out <= 12'h088;
      20'h0bfaf: out <= 12'h088;
      20'h0bfb0: out <= 12'h088;
      20'h0bfb1: out <= 12'h088;
      20'h0bfb2: out <= 12'h088;
      20'h0bfb3: out <= 12'h088;
      20'h0bfb4: out <= 12'h088;
      20'h0bfb5: out <= 12'h088;
      20'h0bfb6: out <= 12'h088;
      20'h0bfb7: out <= 12'h088;
      20'h0bfb8: out <= 12'h088;
      20'h0bfb9: out <= 12'h088;
      20'h0bfba: out <= 12'h088;
      20'h0bfbb: out <= 12'h088;
      20'h0bfbc: out <= 12'h088;
      20'h0bfbd: out <= 12'h088;
      20'h0bfbe: out <= 12'h088;
      20'h0bfbf: out <= 12'h088;
      20'h0bfc0: out <= 12'h088;
      20'h0bfc1: out <= 12'h088;
      20'h0bfc2: out <= 12'h088;
      20'h0bfc3: out <= 12'h088;
      20'h0bfc4: out <= 12'h088;
      20'h0bfc5: out <= 12'h088;
      20'h0bfc6: out <= 12'h088;
      20'h0bfc7: out <= 12'h088;
      20'h0bfc8: out <= 12'h088;
      20'h0bfc9: out <= 12'h088;
      20'h0bfca: out <= 12'h088;
      20'h0bfcb: out <= 12'h088;
      20'h0bfcc: out <= 12'h088;
      20'h0bfcd: out <= 12'h088;
      20'h0bfce: out <= 12'h088;
      20'h0bfcf: out <= 12'h088;
      20'h0bfd0: out <= 12'h088;
      20'h0bfd1: out <= 12'h222;
      20'h0bfd2: out <= 12'h222;
      20'h0bfd3: out <= 12'h660;
      20'h0bfd4: out <= 12'hbb0;
      20'h0bfd5: out <= 12'hee9;
      20'h0bfd6: out <= 12'hee9;
      20'h0bfd7: out <= 12'hee9;
      20'h0bfd8: out <= 12'hee9;
      20'h0bfd9: out <= 12'hee9;
      20'h0bfda: out <= 12'hee9;
      20'h0bfdb: out <= 12'hee9;
      20'h0bfdc: out <= 12'hee9;
      20'h0bfdd: out <= 12'hee9;
      20'h0bfde: out <= 12'hee9;
      20'h0bfdf: out <= 12'hee9;
      20'h0bfe0: out <= 12'hee9;
      20'h0bfe1: out <= 12'hee9;
      20'h0bfe2: out <= 12'hee9;
      20'h0bfe3: out <= 12'hee9;
      20'h0bfe4: out <= 12'hbb0;
      20'h0bfe5: out <= 12'h660;
      20'h0bfe6: out <= 12'h222;
      20'h0bfe7: out <= 12'h222;
      20'h0bfe8: out <= 12'h603;
      20'h0bfe9: out <= 12'h603;
      20'h0bfea: out <= 12'h603;
      20'h0bfeb: out <= 12'h603;
      20'h0bfec: out <= 12'hee9;
      20'h0bfed: out <= 12'hee9;
      20'h0bfee: out <= 12'h000;
      20'h0bfef: out <= 12'hee9;
      20'h0bff0: out <= 12'h000;
      20'h0bff1: out <= 12'hee9;
      20'h0bff2: out <= 12'hee9;
      20'h0bff3: out <= 12'h000;
      20'h0bff4: out <= 12'h000;
      20'h0bff5: out <= 12'h000;
      20'h0bff6: out <= 12'h000;
      20'h0bff7: out <= 12'hee9;
      20'h0bff8: out <= 12'hee9;
      20'h0bff9: out <= 12'h000;
      20'h0bffa: out <= 12'h000;
      20'h0bffb: out <= 12'h000;
      20'h0bffc: out <= 12'h000;
      20'h0bffd: out <= 12'h000;
      20'h0bffe: out <= 12'h000;
      20'h0bfff: out <= 12'hee9;
      20'h0c000: out <= 12'hee9;
      20'h0c001: out <= 12'hee9;
      20'h0c002: out <= 12'h000;
      20'h0c003: out <= 12'h000;
      20'h0c004: out <= 12'h000;
      20'h0c005: out <= 12'h000;
      20'h0c006: out <= 12'hee9;
      20'h0c007: out <= 12'hee9;
      20'h0c008: out <= 12'hee9;
      20'h0c009: out <= 12'hee9;
      20'h0c00a: out <= 12'h000;
      20'h0c00b: out <= 12'h000;
      20'h0c00c: out <= 12'hee9;
      20'h0c00d: out <= 12'hee9;
      20'h0c00e: out <= 12'hee9;
      20'h0c00f: out <= 12'h000;
      20'h0c010: out <= 12'hee9;
      20'h0c011: out <= 12'hee9;
      20'h0c012: out <= 12'h000;
      20'h0c013: out <= 12'h000;
      20'h0c014: out <= 12'h000;
      20'h0c015: out <= 12'h000;
      20'h0c016: out <= 12'h000;
      20'h0c017: out <= 12'h000;
      20'h0c018: out <= 12'h000;
      20'h0c019: out <= 12'hee9;
      20'h0c01a: out <= 12'hee9;
      20'h0c01b: out <= 12'h000;
      20'h0c01c: out <= 12'hee9;
      20'h0c01d: out <= 12'hee9;
      20'h0c01e: out <= 12'hee9;
      20'h0c01f: out <= 12'hee9;
      20'h0c020: out <= 12'hee9;
      20'h0c021: out <= 12'hee9;
      20'h0c022: out <= 12'hee9;
      20'h0c023: out <= 12'h000;
      20'h0c024: out <= 12'h000;
      20'h0c025: out <= 12'h000;
      20'h0c026: out <= 12'h000;
      20'h0c027: out <= 12'hee9;
      20'h0c028: out <= 12'hee9;
      20'h0c029: out <= 12'h000;
      20'h0c02a: out <= 12'h000;
      20'h0c02b: out <= 12'h000;
      20'h0c02c: out <= 12'hee9;
      20'h0c02d: out <= 12'hee9;
      20'h0c02e: out <= 12'hee9;
      20'h0c02f: out <= 12'hee9;
      20'h0c030: out <= 12'hee9;
      20'h0c031: out <= 12'hee9;
      20'h0c032: out <= 12'hee9;
      20'h0c033: out <= 12'h000;
      20'h0c034: out <= 12'h000;
      20'h0c035: out <= 12'hee9;
      20'h0c036: out <= 12'hee9;
      20'h0c037: out <= 12'hee9;
      20'h0c038: out <= 12'hee9;
      20'h0c039: out <= 12'hee9;
      20'h0c03a: out <= 12'hee9;
      20'h0c03b: out <= 12'h000;
      20'h0c03c: out <= 12'h603;
      20'h0c03d: out <= 12'h603;
      20'h0c03e: out <= 12'h603;
      20'h0c03f: out <= 12'h603;
      20'h0c040: out <= 12'hb27;
      20'h0c041: out <= 12'hb27;
      20'h0c042: out <= 12'hb27;
      20'h0c043: out <= 12'hb27;
      20'h0c044: out <= 12'hb27;
      20'h0c045: out <= 12'hb27;
      20'h0c046: out <= 12'hb27;
      20'h0c047: out <= 12'hb27;
      20'h0c048: out <= 12'h000;
      20'h0c049: out <= 12'h000;
      20'h0c04a: out <= 12'h000;
      20'h0c04b: out <= 12'h000;
      20'h0c04c: out <= 12'h000;
      20'h0c04d: out <= 12'h000;
      20'h0c04e: out <= 12'h000;
      20'h0c04f: out <= 12'h000;
      20'h0c050: out <= 12'h777;
      20'h0c051: out <= 12'h777;
      20'h0c052: out <= 12'h777;
      20'h0c053: out <= 12'h777;
      20'h0c054: out <= 12'h777;
      20'h0c055: out <= 12'h777;
      20'h0c056: out <= 12'h777;
      20'h0c057: out <= 12'h777;
      20'h0c058: out <= 12'h777;
      20'h0c059: out <= 12'h777;
      20'h0c05a: out <= 12'h777;
      20'h0c05b: out <= 12'h777;
      20'h0c05c: out <= 12'h777;
      20'h0c05d: out <= 12'h777;
      20'h0c05e: out <= 12'h777;
      20'h0c05f: out <= 12'h777;
      20'h0c060: out <= 12'h000;
      20'h0c061: out <= 12'h000;
      20'h0c062: out <= 12'h000;
      20'h0c063: out <= 12'h000;
      20'h0c064: out <= 12'h000;
      20'h0c065: out <= 12'h000;
      20'h0c066: out <= 12'h000;
      20'h0c067: out <= 12'h000;
      20'h0c068: out <= 12'hfa9;
      20'h0c069: out <= 12'hfa9;
      20'h0c06a: out <= 12'hfa9;
      20'h0c06b: out <= 12'hfa9;
      20'h0c06c: out <= 12'hfa9;
      20'h0c06d: out <= 12'hfa9;
      20'h0c06e: out <= 12'hfa9;
      20'h0c06f: out <= 12'hfa9;
      20'h0c070: out <= 12'hf76;
      20'h0c071: out <= 12'hf76;
      20'h0c072: out <= 12'hf76;
      20'h0c073: out <= 12'hf76;
      20'h0c074: out <= 12'hf76;
      20'h0c075: out <= 12'hf76;
      20'h0c076: out <= 12'hf76;
      20'h0c077: out <= 12'hf76;
      20'h0c078: out <= 12'h000;
      20'h0c079: out <= 12'h000;
      20'h0c07a: out <= 12'h000;
      20'h0c07b: out <= 12'h000;
      20'h0c07c: out <= 12'h000;
      20'h0c07d: out <= 12'h000;
      20'h0c07e: out <= 12'h000;
      20'h0c07f: out <= 12'h000;
      20'h0c080: out <= 12'h088;
      20'h0c081: out <= 12'h088;
      20'h0c082: out <= 12'h088;
      20'h0c083: out <= 12'h088;
      20'h0c084: out <= 12'h088;
      20'h0c085: out <= 12'h088;
      20'h0c086: out <= 12'h088;
      20'h0c087: out <= 12'h088;
      20'h0c088: out <= 12'h088;
      20'h0c089: out <= 12'h088;
      20'h0c08a: out <= 12'h088;
      20'h0c08b: out <= 12'h088;
      20'h0c08c: out <= 12'h088;
      20'h0c08d: out <= 12'h088;
      20'h0c08e: out <= 12'h088;
      20'h0c08f: out <= 12'h088;
      20'h0c090: out <= 12'h088;
      20'h0c091: out <= 12'h088;
      20'h0c092: out <= 12'h088;
      20'h0c093: out <= 12'h088;
      20'h0c094: out <= 12'h088;
      20'h0c095: out <= 12'h088;
      20'h0c096: out <= 12'h088;
      20'h0c097: out <= 12'h088;
      20'h0c098: out <= 12'h088;
      20'h0c099: out <= 12'h088;
      20'h0c09a: out <= 12'h088;
      20'h0c09b: out <= 12'h088;
      20'h0c09c: out <= 12'h088;
      20'h0c09d: out <= 12'h088;
      20'h0c09e: out <= 12'h088;
      20'h0c09f: out <= 12'h088;
      20'h0c0a0: out <= 12'h088;
      20'h0c0a1: out <= 12'h088;
      20'h0c0a2: out <= 12'h088;
      20'h0c0a3: out <= 12'h088;
      20'h0c0a4: out <= 12'h088;
      20'h0c0a5: out <= 12'h088;
      20'h0c0a6: out <= 12'h088;
      20'h0c0a7: out <= 12'h088;
      20'h0c0a8: out <= 12'h088;
      20'h0c0a9: out <= 12'h088;
      20'h0c0aa: out <= 12'h088;
      20'h0c0ab: out <= 12'h088;
      20'h0c0ac: out <= 12'h088;
      20'h0c0ad: out <= 12'h088;
      20'h0c0ae: out <= 12'h088;
      20'h0c0af: out <= 12'h088;
      20'h0c0b0: out <= 12'h088;
      20'h0c0b1: out <= 12'h088;
      20'h0c0b2: out <= 12'h088;
      20'h0c0b3: out <= 12'h088;
      20'h0c0b4: out <= 12'h088;
      20'h0c0b5: out <= 12'h088;
      20'h0c0b6: out <= 12'h088;
      20'h0c0b7: out <= 12'h088;
      20'h0c0b8: out <= 12'h088;
      20'h0c0b9: out <= 12'h088;
      20'h0c0ba: out <= 12'h088;
      20'h0c0bb: out <= 12'h088;
      20'h0c0bc: out <= 12'h088;
      20'h0c0bd: out <= 12'h088;
      20'h0c0be: out <= 12'h088;
      20'h0c0bf: out <= 12'h088;
      20'h0c0c0: out <= 12'h088;
      20'h0c0c1: out <= 12'h088;
      20'h0c0c2: out <= 12'h088;
      20'h0c0c3: out <= 12'h088;
      20'h0c0c4: out <= 12'h088;
      20'h0c0c5: out <= 12'h088;
      20'h0c0c6: out <= 12'h088;
      20'h0c0c7: out <= 12'h088;
      20'h0c0c8: out <= 12'h088;
      20'h0c0c9: out <= 12'h088;
      20'h0c0ca: out <= 12'h088;
      20'h0c0cb: out <= 12'h088;
      20'h0c0cc: out <= 12'h088;
      20'h0c0cd: out <= 12'h088;
      20'h0c0ce: out <= 12'h088;
      20'h0c0cf: out <= 12'h088;
      20'h0c0d0: out <= 12'h088;
      20'h0c0d1: out <= 12'h088;
      20'h0c0d2: out <= 12'h088;
      20'h0c0d3: out <= 12'h088;
      20'h0c0d4: out <= 12'h088;
      20'h0c0d5: out <= 12'h088;
      20'h0c0d6: out <= 12'h088;
      20'h0c0d7: out <= 12'h088;
      20'h0c0d8: out <= 12'h088;
      20'h0c0d9: out <= 12'h088;
      20'h0c0da: out <= 12'h088;
      20'h0c0db: out <= 12'h088;
      20'h0c0dc: out <= 12'h088;
      20'h0c0dd: out <= 12'h088;
      20'h0c0de: out <= 12'h088;
      20'h0c0df: out <= 12'h088;
      20'h0c0e0: out <= 12'h088;
      20'h0c0e1: out <= 12'h088;
      20'h0c0e2: out <= 12'h088;
      20'h0c0e3: out <= 12'h088;
      20'h0c0e4: out <= 12'h088;
      20'h0c0e5: out <= 12'h088;
      20'h0c0e6: out <= 12'h088;
      20'h0c0e7: out <= 12'h088;
      20'h0c0e8: out <= 12'h088;
      20'h0c0e9: out <= 12'h222;
      20'h0c0ea: out <= 12'h222;
      20'h0c0eb: out <= 12'h222;
      20'h0c0ec: out <= 12'h222;
      20'h0c0ed: out <= 12'h660;
      20'h0c0ee: out <= 12'hbb0;
      20'h0c0ef: out <= 12'hee9;
      20'h0c0f0: out <= 12'hee9;
      20'h0c0f1: out <= 12'hee9;
      20'h0c0f2: out <= 12'hee9;
      20'h0c0f3: out <= 12'hee9;
      20'h0c0f4: out <= 12'hee9;
      20'h0c0f5: out <= 12'hee9;
      20'h0c0f6: out <= 12'hee9;
      20'h0c0f7: out <= 12'hee9;
      20'h0c0f8: out <= 12'hee9;
      20'h0c0f9: out <= 12'hee9;
      20'h0c0fa: out <= 12'hbb0;
      20'h0c0fb: out <= 12'h660;
      20'h0c0fc: out <= 12'h222;
      20'h0c0fd: out <= 12'h222;
      20'h0c0fe: out <= 12'h222;
      20'h0c0ff: out <= 12'h222;
      20'h0c100: out <= 12'h603;
      20'h0c101: out <= 12'h603;
      20'h0c102: out <= 12'h603;
      20'h0c103: out <= 12'h603;
      20'h0c104: out <= 12'hee9;
      20'h0c105: out <= 12'hee9;
      20'h0c106: out <= 12'hee9;
      20'h0c107: out <= 12'h000;
      20'h0c108: out <= 12'h000;
      20'h0c109: out <= 12'hee9;
      20'h0c10a: out <= 12'hee9;
      20'h0c10b: out <= 12'h000;
      20'h0c10c: out <= 12'h000;
      20'h0c10d: out <= 12'h000;
      20'h0c10e: out <= 12'h000;
      20'h0c10f: out <= 12'hee9;
      20'h0c110: out <= 12'hee9;
      20'h0c111: out <= 12'h000;
      20'h0c112: out <= 12'h000;
      20'h0c113: out <= 12'h000;
      20'h0c114: out <= 12'h000;
      20'h0c115: out <= 12'h000;
      20'h0c116: out <= 12'hee9;
      20'h0c117: out <= 12'hee9;
      20'h0c118: out <= 12'hee9;
      20'h0c119: out <= 12'h000;
      20'h0c11a: out <= 12'h000;
      20'h0c11b: out <= 12'h000;
      20'h0c11c: out <= 12'h000;
      20'h0c11d: out <= 12'h000;
      20'h0c11e: out <= 12'h000;
      20'h0c11f: out <= 12'h000;
      20'h0c120: out <= 12'h000;
      20'h0c121: out <= 12'hee9;
      20'h0c122: out <= 12'hee9;
      20'h0c123: out <= 12'h000;
      20'h0c124: out <= 12'hee9;
      20'h0c125: out <= 12'hee9;
      20'h0c126: out <= 12'h000;
      20'h0c127: out <= 12'h000;
      20'h0c128: out <= 12'hee9;
      20'h0c129: out <= 12'hee9;
      20'h0c12a: out <= 12'h000;
      20'h0c12b: out <= 12'h000;
      20'h0c12c: out <= 12'h000;
      20'h0c12d: out <= 12'h000;
      20'h0c12e: out <= 12'h000;
      20'h0c12f: out <= 12'h000;
      20'h0c130: out <= 12'h000;
      20'h0c131: out <= 12'hee9;
      20'h0c132: out <= 12'hee9;
      20'h0c133: out <= 12'h000;
      20'h0c134: out <= 12'hee9;
      20'h0c135: out <= 12'hee9;
      20'h0c136: out <= 12'h000;
      20'h0c137: out <= 12'h000;
      20'h0c138: out <= 12'h000;
      20'h0c139: out <= 12'hee9;
      20'h0c13a: out <= 12'hee9;
      20'h0c13b: out <= 12'h000;
      20'h0c13c: out <= 12'h000;
      20'h0c13d: out <= 12'h000;
      20'h0c13e: out <= 12'h000;
      20'h0c13f: out <= 12'hee9;
      20'h0c140: out <= 12'hee9;
      20'h0c141: out <= 12'h000;
      20'h0c142: out <= 12'h000;
      20'h0c143: out <= 12'h000;
      20'h0c144: out <= 12'hee9;
      20'h0c145: out <= 12'hee9;
      20'h0c146: out <= 12'h000;
      20'h0c147: out <= 12'h000;
      20'h0c148: out <= 12'h000;
      20'h0c149: out <= 12'hee9;
      20'h0c14a: out <= 12'hee9;
      20'h0c14b: out <= 12'h000;
      20'h0c14c: out <= 12'h000;
      20'h0c14d: out <= 12'h000;
      20'h0c14e: out <= 12'h000;
      20'h0c14f: out <= 12'h000;
      20'h0c150: out <= 12'h000;
      20'h0c151: out <= 12'hee9;
      20'h0c152: out <= 12'hee9;
      20'h0c153: out <= 12'h000;
      20'h0c154: out <= 12'h603;
      20'h0c155: out <= 12'h603;
      20'h0c156: out <= 12'h603;
      20'h0c157: out <= 12'h603;
      20'h0c158: out <= 12'hee9;
      20'h0c159: out <= 12'hee9;
      20'h0c15a: out <= 12'hee9;
      20'h0c15b: out <= 12'hee9;
      20'h0c15c: out <= 12'hee9;
      20'h0c15d: out <= 12'hee9;
      20'h0c15e: out <= 12'hee9;
      20'h0c15f: out <= 12'hb27;
      20'h0c160: out <= 12'hee9;
      20'h0c161: out <= 12'hee9;
      20'h0c162: out <= 12'hee9;
      20'h0c163: out <= 12'hee9;
      20'h0c164: out <= 12'hee9;
      20'h0c165: out <= 12'hee9;
      20'h0c166: out <= 12'hee9;
      20'h0c167: out <= 12'hb27;
      20'h0c168: out <= 12'hee9;
      20'h0c169: out <= 12'hee9;
      20'h0c16a: out <= 12'hee9;
      20'h0c16b: out <= 12'hee9;
      20'h0c16c: out <= 12'hee9;
      20'h0c16d: out <= 12'hee9;
      20'h0c16e: out <= 12'hee9;
      20'h0c16f: out <= 12'hb27;
      20'h0c170: out <= 12'hee9;
      20'h0c171: out <= 12'hee9;
      20'h0c172: out <= 12'hee9;
      20'h0c173: out <= 12'hee9;
      20'h0c174: out <= 12'hee9;
      20'h0c175: out <= 12'hee9;
      20'h0c176: out <= 12'hee9;
      20'h0c177: out <= 12'hb27;
      20'h0c178: out <= 12'hee9;
      20'h0c179: out <= 12'hee9;
      20'h0c17a: out <= 12'hee9;
      20'h0c17b: out <= 12'hee9;
      20'h0c17c: out <= 12'hee9;
      20'h0c17d: out <= 12'hee9;
      20'h0c17e: out <= 12'hee9;
      20'h0c17f: out <= 12'hb27;
      20'h0c180: out <= 12'hee9;
      20'h0c181: out <= 12'hee9;
      20'h0c182: out <= 12'hee9;
      20'h0c183: out <= 12'hee9;
      20'h0c184: out <= 12'hee9;
      20'h0c185: out <= 12'hee9;
      20'h0c186: out <= 12'hee9;
      20'h0c187: out <= 12'hb27;
      20'h0c188: out <= 12'hee9;
      20'h0c189: out <= 12'hee9;
      20'h0c18a: out <= 12'hee9;
      20'h0c18b: out <= 12'hee9;
      20'h0c18c: out <= 12'hee9;
      20'h0c18d: out <= 12'hee9;
      20'h0c18e: out <= 12'hee9;
      20'h0c18f: out <= 12'hb27;
      20'h0c190: out <= 12'hee9;
      20'h0c191: out <= 12'hee9;
      20'h0c192: out <= 12'hee9;
      20'h0c193: out <= 12'hee9;
      20'h0c194: out <= 12'hee9;
      20'h0c195: out <= 12'hee9;
      20'h0c196: out <= 12'hee9;
      20'h0c197: out <= 12'hb27;
      20'h0c198: out <= 12'h088;
      20'h0c199: out <= 12'h088;
      20'h0c19a: out <= 12'h088;
      20'h0c19b: out <= 12'h088;
      20'h0c19c: out <= 12'h088;
      20'h0c19d: out <= 12'h088;
      20'h0c19e: out <= 12'h088;
      20'h0c19f: out <= 12'h088;
      20'h0c1a0: out <= 12'h088;
      20'h0c1a1: out <= 12'h088;
      20'h0c1a2: out <= 12'h088;
      20'h0c1a3: out <= 12'h088;
      20'h0c1a4: out <= 12'h088;
      20'h0c1a5: out <= 12'h088;
      20'h0c1a6: out <= 12'h088;
      20'h0c1a7: out <= 12'h088;
      20'h0c1a8: out <= 12'h088;
      20'h0c1a9: out <= 12'h088;
      20'h0c1aa: out <= 12'h088;
      20'h0c1ab: out <= 12'h088;
      20'h0c1ac: out <= 12'h088;
      20'h0c1ad: out <= 12'h088;
      20'h0c1ae: out <= 12'h088;
      20'h0c1af: out <= 12'h088;
      20'h0c1b0: out <= 12'h088;
      20'h0c1b1: out <= 12'h088;
      20'h0c1b2: out <= 12'h088;
      20'h0c1b3: out <= 12'h088;
      20'h0c1b4: out <= 12'h088;
      20'h0c1b5: out <= 12'h088;
      20'h0c1b6: out <= 12'h088;
      20'h0c1b7: out <= 12'h088;
      20'h0c1b8: out <= 12'h088;
      20'h0c1b9: out <= 12'h088;
      20'h0c1ba: out <= 12'h088;
      20'h0c1bb: out <= 12'h088;
      20'h0c1bc: out <= 12'h088;
      20'h0c1bd: out <= 12'h088;
      20'h0c1be: out <= 12'h088;
      20'h0c1bf: out <= 12'h088;
      20'h0c1c0: out <= 12'h088;
      20'h0c1c1: out <= 12'h088;
      20'h0c1c2: out <= 12'h088;
      20'h0c1c3: out <= 12'h088;
      20'h0c1c4: out <= 12'h088;
      20'h0c1c5: out <= 12'h088;
      20'h0c1c6: out <= 12'h088;
      20'h0c1c7: out <= 12'h088;
      20'h0c1c8: out <= 12'h088;
      20'h0c1c9: out <= 12'h088;
      20'h0c1ca: out <= 12'h088;
      20'h0c1cb: out <= 12'h088;
      20'h0c1cc: out <= 12'h088;
      20'h0c1cd: out <= 12'h088;
      20'h0c1ce: out <= 12'h088;
      20'h0c1cf: out <= 12'h088;
      20'h0c1d0: out <= 12'h088;
      20'h0c1d1: out <= 12'h088;
      20'h0c1d2: out <= 12'h088;
      20'h0c1d3: out <= 12'h088;
      20'h0c1d4: out <= 12'h088;
      20'h0c1d5: out <= 12'h088;
      20'h0c1d6: out <= 12'h088;
      20'h0c1d7: out <= 12'h088;
      20'h0c1d8: out <= 12'h088;
      20'h0c1d9: out <= 12'h088;
      20'h0c1da: out <= 12'h088;
      20'h0c1db: out <= 12'h088;
      20'h0c1dc: out <= 12'h088;
      20'h0c1dd: out <= 12'h088;
      20'h0c1de: out <= 12'h088;
      20'h0c1df: out <= 12'h088;
      20'h0c1e0: out <= 12'h088;
      20'h0c1e1: out <= 12'h088;
      20'h0c1e2: out <= 12'h088;
      20'h0c1e3: out <= 12'h088;
      20'h0c1e4: out <= 12'h088;
      20'h0c1e5: out <= 12'h088;
      20'h0c1e6: out <= 12'h088;
      20'h0c1e7: out <= 12'h088;
      20'h0c1e8: out <= 12'h088;
      20'h0c1e9: out <= 12'h088;
      20'h0c1ea: out <= 12'h088;
      20'h0c1eb: out <= 12'h088;
      20'h0c1ec: out <= 12'h088;
      20'h0c1ed: out <= 12'h088;
      20'h0c1ee: out <= 12'h088;
      20'h0c1ef: out <= 12'h088;
      20'h0c1f0: out <= 12'h088;
      20'h0c1f1: out <= 12'h088;
      20'h0c1f2: out <= 12'h088;
      20'h0c1f3: out <= 12'h088;
      20'h0c1f4: out <= 12'h088;
      20'h0c1f5: out <= 12'h088;
      20'h0c1f6: out <= 12'h088;
      20'h0c1f7: out <= 12'h088;
      20'h0c1f8: out <= 12'h088;
      20'h0c1f9: out <= 12'h088;
      20'h0c1fa: out <= 12'h088;
      20'h0c1fb: out <= 12'h088;
      20'h0c1fc: out <= 12'h088;
      20'h0c1fd: out <= 12'h088;
      20'h0c1fe: out <= 12'h088;
      20'h0c1ff: out <= 12'h088;
      20'h0c200: out <= 12'h088;
      20'h0c201: out <= 12'h222;
      20'h0c202: out <= 12'h222;
      20'h0c203: out <= 12'h222;
      20'h0c204: out <= 12'h222;
      20'h0c205: out <= 12'h222;
      20'h0c206: out <= 12'h660;
      20'h0c207: out <= 12'hbb0;
      20'h0c208: out <= 12'hee9;
      20'h0c209: out <= 12'hee9;
      20'h0c20a: out <= 12'hee9;
      20'h0c20b: out <= 12'hee9;
      20'h0c20c: out <= 12'hee9;
      20'h0c20d: out <= 12'hee9;
      20'h0c20e: out <= 12'hee9;
      20'h0c20f: out <= 12'hee9;
      20'h0c210: out <= 12'hee9;
      20'h0c211: out <= 12'hbb0;
      20'h0c212: out <= 12'h660;
      20'h0c213: out <= 12'h222;
      20'h0c214: out <= 12'h222;
      20'h0c215: out <= 12'h222;
      20'h0c216: out <= 12'h222;
      20'h0c217: out <= 12'h222;
      20'h0c218: out <= 12'h603;
      20'h0c219: out <= 12'h603;
      20'h0c21a: out <= 12'h603;
      20'h0c21b: out <= 12'h603;
      20'h0c21c: out <= 12'hee9;
      20'h0c21d: out <= 12'hee9;
      20'h0c21e: out <= 12'hee9;
      20'h0c21f: out <= 12'h000;
      20'h0c220: out <= 12'h000;
      20'h0c221: out <= 12'hee9;
      20'h0c222: out <= 12'hee9;
      20'h0c223: out <= 12'h000;
      20'h0c224: out <= 12'h000;
      20'h0c225: out <= 12'h000;
      20'h0c226: out <= 12'h000;
      20'h0c227: out <= 12'hee9;
      20'h0c228: out <= 12'hee9;
      20'h0c229: out <= 12'h000;
      20'h0c22a: out <= 12'h000;
      20'h0c22b: out <= 12'h000;
      20'h0c22c: out <= 12'h000;
      20'h0c22d: out <= 12'hee9;
      20'h0c22e: out <= 12'hee9;
      20'h0c22f: out <= 12'hee9;
      20'h0c230: out <= 12'h000;
      20'h0c231: out <= 12'h000;
      20'h0c232: out <= 12'h000;
      20'h0c233: out <= 12'h000;
      20'h0c234: out <= 12'h000;
      20'h0c235: out <= 12'h000;
      20'h0c236: out <= 12'h000;
      20'h0c237: out <= 12'h000;
      20'h0c238: out <= 12'h000;
      20'h0c239: out <= 12'hee9;
      20'h0c23a: out <= 12'hee9;
      20'h0c23b: out <= 12'h000;
      20'h0c23c: out <= 12'hee9;
      20'h0c23d: out <= 12'hee9;
      20'h0c23e: out <= 12'h000;
      20'h0c23f: out <= 12'h000;
      20'h0c240: out <= 12'hee9;
      20'h0c241: out <= 12'hee9;
      20'h0c242: out <= 12'h000;
      20'h0c243: out <= 12'h000;
      20'h0c244: out <= 12'h000;
      20'h0c245: out <= 12'h000;
      20'h0c246: out <= 12'h000;
      20'h0c247: out <= 12'h000;
      20'h0c248: out <= 12'h000;
      20'h0c249: out <= 12'hee9;
      20'h0c24a: out <= 12'hee9;
      20'h0c24b: out <= 12'h000;
      20'h0c24c: out <= 12'hee9;
      20'h0c24d: out <= 12'hee9;
      20'h0c24e: out <= 12'h000;
      20'h0c24f: out <= 12'h000;
      20'h0c250: out <= 12'h000;
      20'h0c251: out <= 12'hee9;
      20'h0c252: out <= 12'hee9;
      20'h0c253: out <= 12'h000;
      20'h0c254: out <= 12'h000;
      20'h0c255: out <= 12'h000;
      20'h0c256: out <= 12'hee9;
      20'h0c257: out <= 12'hee9;
      20'h0c258: out <= 12'h000;
      20'h0c259: out <= 12'h000;
      20'h0c25a: out <= 12'h000;
      20'h0c25b: out <= 12'h000;
      20'h0c25c: out <= 12'hee9;
      20'h0c25d: out <= 12'hee9;
      20'h0c25e: out <= 12'h000;
      20'h0c25f: out <= 12'h000;
      20'h0c260: out <= 12'h000;
      20'h0c261: out <= 12'hee9;
      20'h0c262: out <= 12'hee9;
      20'h0c263: out <= 12'h000;
      20'h0c264: out <= 12'h000;
      20'h0c265: out <= 12'h000;
      20'h0c266: out <= 12'h000;
      20'h0c267: out <= 12'h000;
      20'h0c268: out <= 12'hee9;
      20'h0c269: out <= 12'hee9;
      20'h0c26a: out <= 12'hee9;
      20'h0c26b: out <= 12'h000;
      20'h0c26c: out <= 12'h603;
      20'h0c26d: out <= 12'h603;
      20'h0c26e: out <= 12'h603;
      20'h0c26f: out <= 12'h603;
      20'h0c270: out <= 12'hee9;
      20'h0c271: out <= 12'hf87;
      20'h0c272: out <= 12'hf87;
      20'h0c273: out <= 12'hf87;
      20'h0c274: out <= 12'hf87;
      20'h0c275: out <= 12'hf87;
      20'h0c276: out <= 12'hf87;
      20'h0c277: out <= 12'hb27;
      20'h0c278: out <= 12'hee9;
      20'h0c279: out <= 12'hf87;
      20'h0c27a: out <= 12'hf87;
      20'h0c27b: out <= 12'hf87;
      20'h0c27c: out <= 12'hf87;
      20'h0c27d: out <= 12'hf87;
      20'h0c27e: out <= 12'hf87;
      20'h0c27f: out <= 12'hb27;
      20'h0c280: out <= 12'hee9;
      20'h0c281: out <= 12'hf87;
      20'h0c282: out <= 12'hf87;
      20'h0c283: out <= 12'hf87;
      20'h0c284: out <= 12'hf87;
      20'h0c285: out <= 12'hf87;
      20'h0c286: out <= 12'hf87;
      20'h0c287: out <= 12'hb27;
      20'h0c288: out <= 12'hee9;
      20'h0c289: out <= 12'hf87;
      20'h0c28a: out <= 12'hf87;
      20'h0c28b: out <= 12'hf87;
      20'h0c28c: out <= 12'hf87;
      20'h0c28d: out <= 12'hf87;
      20'h0c28e: out <= 12'hf87;
      20'h0c28f: out <= 12'hb27;
      20'h0c290: out <= 12'hee9;
      20'h0c291: out <= 12'hf87;
      20'h0c292: out <= 12'hf87;
      20'h0c293: out <= 12'hf87;
      20'h0c294: out <= 12'hf87;
      20'h0c295: out <= 12'hf87;
      20'h0c296: out <= 12'hf87;
      20'h0c297: out <= 12'hb27;
      20'h0c298: out <= 12'hee9;
      20'h0c299: out <= 12'hf87;
      20'h0c29a: out <= 12'hf87;
      20'h0c29b: out <= 12'hf87;
      20'h0c29c: out <= 12'hf87;
      20'h0c29d: out <= 12'hf87;
      20'h0c29e: out <= 12'hf87;
      20'h0c29f: out <= 12'hb27;
      20'h0c2a0: out <= 12'hee9;
      20'h0c2a1: out <= 12'hf87;
      20'h0c2a2: out <= 12'hf87;
      20'h0c2a3: out <= 12'hf87;
      20'h0c2a4: out <= 12'hf87;
      20'h0c2a5: out <= 12'hf87;
      20'h0c2a6: out <= 12'hf87;
      20'h0c2a7: out <= 12'hb27;
      20'h0c2a8: out <= 12'hee9;
      20'h0c2a9: out <= 12'hf87;
      20'h0c2aa: out <= 12'hf87;
      20'h0c2ab: out <= 12'hf87;
      20'h0c2ac: out <= 12'hf87;
      20'h0c2ad: out <= 12'hf87;
      20'h0c2ae: out <= 12'hf87;
      20'h0c2af: out <= 12'hb27;
      20'h0c2b0: out <= 12'h088;
      20'h0c2b1: out <= 12'h088;
      20'h0c2b2: out <= 12'h088;
      20'h0c2b3: out <= 12'h088;
      20'h0c2b4: out <= 12'h088;
      20'h0c2b5: out <= 12'h088;
      20'h0c2b6: out <= 12'h088;
      20'h0c2b7: out <= 12'h088;
      20'h0c2b8: out <= 12'h088;
      20'h0c2b9: out <= 12'h088;
      20'h0c2ba: out <= 12'h088;
      20'h0c2bb: out <= 12'h088;
      20'h0c2bc: out <= 12'h088;
      20'h0c2bd: out <= 12'h088;
      20'h0c2be: out <= 12'h088;
      20'h0c2bf: out <= 12'h088;
      20'h0c2c0: out <= 12'h088;
      20'h0c2c1: out <= 12'h088;
      20'h0c2c2: out <= 12'h088;
      20'h0c2c3: out <= 12'h088;
      20'h0c2c4: out <= 12'h088;
      20'h0c2c5: out <= 12'h088;
      20'h0c2c6: out <= 12'h088;
      20'h0c2c7: out <= 12'h088;
      20'h0c2c8: out <= 12'h088;
      20'h0c2c9: out <= 12'h088;
      20'h0c2ca: out <= 12'h088;
      20'h0c2cb: out <= 12'h088;
      20'h0c2cc: out <= 12'h088;
      20'h0c2cd: out <= 12'h088;
      20'h0c2ce: out <= 12'h088;
      20'h0c2cf: out <= 12'h088;
      20'h0c2d0: out <= 12'h088;
      20'h0c2d1: out <= 12'h088;
      20'h0c2d2: out <= 12'h088;
      20'h0c2d3: out <= 12'h088;
      20'h0c2d4: out <= 12'h088;
      20'h0c2d5: out <= 12'h088;
      20'h0c2d6: out <= 12'h088;
      20'h0c2d7: out <= 12'h088;
      20'h0c2d8: out <= 12'h088;
      20'h0c2d9: out <= 12'h088;
      20'h0c2da: out <= 12'h088;
      20'h0c2db: out <= 12'h088;
      20'h0c2dc: out <= 12'h088;
      20'h0c2dd: out <= 12'h088;
      20'h0c2de: out <= 12'h088;
      20'h0c2df: out <= 12'h088;
      20'h0c2e0: out <= 12'h088;
      20'h0c2e1: out <= 12'h088;
      20'h0c2e2: out <= 12'h088;
      20'h0c2e3: out <= 12'h088;
      20'h0c2e4: out <= 12'h088;
      20'h0c2e5: out <= 12'h088;
      20'h0c2e6: out <= 12'h088;
      20'h0c2e7: out <= 12'h088;
      20'h0c2e8: out <= 12'h088;
      20'h0c2e9: out <= 12'h088;
      20'h0c2ea: out <= 12'h088;
      20'h0c2eb: out <= 12'h088;
      20'h0c2ec: out <= 12'h088;
      20'h0c2ed: out <= 12'h088;
      20'h0c2ee: out <= 12'h088;
      20'h0c2ef: out <= 12'h088;
      20'h0c2f0: out <= 12'h088;
      20'h0c2f1: out <= 12'h088;
      20'h0c2f2: out <= 12'h088;
      20'h0c2f3: out <= 12'h088;
      20'h0c2f4: out <= 12'h088;
      20'h0c2f5: out <= 12'h088;
      20'h0c2f6: out <= 12'h088;
      20'h0c2f7: out <= 12'h088;
      20'h0c2f8: out <= 12'h088;
      20'h0c2f9: out <= 12'h088;
      20'h0c2fa: out <= 12'h088;
      20'h0c2fb: out <= 12'h088;
      20'h0c2fc: out <= 12'h088;
      20'h0c2fd: out <= 12'h088;
      20'h0c2fe: out <= 12'h088;
      20'h0c2ff: out <= 12'h088;
      20'h0c300: out <= 12'h088;
      20'h0c301: out <= 12'h088;
      20'h0c302: out <= 12'h088;
      20'h0c303: out <= 12'h088;
      20'h0c304: out <= 12'h088;
      20'h0c305: out <= 12'h088;
      20'h0c306: out <= 12'h088;
      20'h0c307: out <= 12'h088;
      20'h0c308: out <= 12'h088;
      20'h0c309: out <= 12'h088;
      20'h0c30a: out <= 12'h088;
      20'h0c30b: out <= 12'h088;
      20'h0c30c: out <= 12'h088;
      20'h0c30d: out <= 12'h088;
      20'h0c30e: out <= 12'h088;
      20'h0c30f: out <= 12'h088;
      20'h0c310: out <= 12'h088;
      20'h0c311: out <= 12'h088;
      20'h0c312: out <= 12'h088;
      20'h0c313: out <= 12'h088;
      20'h0c314: out <= 12'h088;
      20'h0c315: out <= 12'h088;
      20'h0c316: out <= 12'h088;
      20'h0c317: out <= 12'h088;
      20'h0c318: out <= 12'h088;
      20'h0c319: out <= 12'h222;
      20'h0c31a: out <= 12'h222;
      20'h0c31b: out <= 12'h222;
      20'h0c31c: out <= 12'h222;
      20'h0c31d: out <= 12'h222;
      20'h0c31e: out <= 12'h222;
      20'h0c31f: out <= 12'h660;
      20'h0c320: out <= 12'hbb0;
      20'h0c321: out <= 12'hee9;
      20'h0c322: out <= 12'hee9;
      20'h0c323: out <= 12'hee9;
      20'h0c324: out <= 12'hee9;
      20'h0c325: out <= 12'hee9;
      20'h0c326: out <= 12'hee9;
      20'h0c327: out <= 12'hee9;
      20'h0c328: out <= 12'hbb0;
      20'h0c329: out <= 12'h660;
      20'h0c32a: out <= 12'h222;
      20'h0c32b: out <= 12'h222;
      20'h0c32c: out <= 12'h222;
      20'h0c32d: out <= 12'h222;
      20'h0c32e: out <= 12'h222;
      20'h0c32f: out <= 12'h222;
      20'h0c330: out <= 12'h603;
      20'h0c331: out <= 12'h603;
      20'h0c332: out <= 12'h603;
      20'h0c333: out <= 12'h603;
      20'h0c334: out <= 12'hf87;
      20'h0c335: out <= 12'hf87;
      20'h0c336: out <= 12'h000;
      20'h0c337: out <= 12'h000;
      20'h0c338: out <= 12'h000;
      20'h0c339: out <= 12'hf87;
      20'h0c33a: out <= 12'hf87;
      20'h0c33b: out <= 12'h000;
      20'h0c33c: out <= 12'h000;
      20'h0c33d: out <= 12'h000;
      20'h0c33e: out <= 12'h000;
      20'h0c33f: out <= 12'hf87;
      20'h0c340: out <= 12'hf87;
      20'h0c341: out <= 12'h000;
      20'h0c342: out <= 12'h000;
      20'h0c343: out <= 12'h000;
      20'h0c344: out <= 12'h000;
      20'h0c345: out <= 12'hf87;
      20'h0c346: out <= 12'hf87;
      20'h0c347: out <= 12'h000;
      20'h0c348: out <= 12'h000;
      20'h0c349: out <= 12'h000;
      20'h0c34a: out <= 12'h000;
      20'h0c34b: out <= 12'h000;
      20'h0c34c: out <= 12'hf87;
      20'h0c34d: out <= 12'hf87;
      20'h0c34e: out <= 12'h000;
      20'h0c34f: out <= 12'h000;
      20'h0c350: out <= 12'h000;
      20'h0c351: out <= 12'hf87;
      20'h0c352: out <= 12'hf87;
      20'h0c353: out <= 12'h000;
      20'h0c354: out <= 12'hf87;
      20'h0c355: out <= 12'hf87;
      20'h0c356: out <= 12'hf87;
      20'h0c357: out <= 12'hf87;
      20'h0c358: out <= 12'hf87;
      20'h0c359: out <= 12'hf87;
      20'h0c35a: out <= 12'hf87;
      20'h0c35b: out <= 12'h000;
      20'h0c35c: out <= 12'hf87;
      20'h0c35d: out <= 12'hf87;
      20'h0c35e: out <= 12'h000;
      20'h0c35f: out <= 12'h000;
      20'h0c360: out <= 12'h000;
      20'h0c361: out <= 12'hf87;
      20'h0c362: out <= 12'hf87;
      20'h0c363: out <= 12'h000;
      20'h0c364: out <= 12'hf87;
      20'h0c365: out <= 12'hf87;
      20'h0c366: out <= 12'h000;
      20'h0c367: out <= 12'h000;
      20'h0c368: out <= 12'h000;
      20'h0c369: out <= 12'hf87;
      20'h0c36a: out <= 12'hf87;
      20'h0c36b: out <= 12'h000;
      20'h0c36c: out <= 12'h000;
      20'h0c36d: out <= 12'h000;
      20'h0c36e: out <= 12'hf87;
      20'h0c36f: out <= 12'hf87;
      20'h0c370: out <= 12'h000;
      20'h0c371: out <= 12'h000;
      20'h0c372: out <= 12'h000;
      20'h0c373: out <= 12'h000;
      20'h0c374: out <= 12'hf87;
      20'h0c375: out <= 12'hf87;
      20'h0c376: out <= 12'h000;
      20'h0c377: out <= 12'h000;
      20'h0c378: out <= 12'h000;
      20'h0c379: out <= 12'hf87;
      20'h0c37a: out <= 12'hf87;
      20'h0c37b: out <= 12'h000;
      20'h0c37c: out <= 12'h000;
      20'h0c37d: out <= 12'h000;
      20'h0c37e: out <= 12'h000;
      20'h0c37f: out <= 12'h000;
      20'h0c380: out <= 12'hf87;
      20'h0c381: out <= 12'hf87;
      20'h0c382: out <= 12'h000;
      20'h0c383: out <= 12'h000;
      20'h0c384: out <= 12'h603;
      20'h0c385: out <= 12'h603;
      20'h0c386: out <= 12'h603;
      20'h0c387: out <= 12'h603;
      20'h0c388: out <= 12'hee9;
      20'h0c389: out <= 12'hf87;
      20'h0c38a: out <= 12'hee9;
      20'h0c38b: out <= 12'hee9;
      20'h0c38c: out <= 12'hee9;
      20'h0c38d: out <= 12'hb27;
      20'h0c38e: out <= 12'hf87;
      20'h0c38f: out <= 12'hb27;
      20'h0c390: out <= 12'hee9;
      20'h0c391: out <= 12'hf87;
      20'h0c392: out <= 12'hee9;
      20'h0c393: out <= 12'hee9;
      20'h0c394: out <= 12'hee9;
      20'h0c395: out <= 12'hb27;
      20'h0c396: out <= 12'hf87;
      20'h0c397: out <= 12'hb27;
      20'h0c398: out <= 12'hee9;
      20'h0c399: out <= 12'hf87;
      20'h0c39a: out <= 12'hee9;
      20'h0c39b: out <= 12'hee9;
      20'h0c39c: out <= 12'hee9;
      20'h0c39d: out <= 12'hb27;
      20'h0c39e: out <= 12'hf87;
      20'h0c39f: out <= 12'hb27;
      20'h0c3a0: out <= 12'hee9;
      20'h0c3a1: out <= 12'hf87;
      20'h0c3a2: out <= 12'hee9;
      20'h0c3a3: out <= 12'hee9;
      20'h0c3a4: out <= 12'hee9;
      20'h0c3a5: out <= 12'hb27;
      20'h0c3a6: out <= 12'hf87;
      20'h0c3a7: out <= 12'hb27;
      20'h0c3a8: out <= 12'hee9;
      20'h0c3a9: out <= 12'hf87;
      20'h0c3aa: out <= 12'hee9;
      20'h0c3ab: out <= 12'hee9;
      20'h0c3ac: out <= 12'hee9;
      20'h0c3ad: out <= 12'hb27;
      20'h0c3ae: out <= 12'hf87;
      20'h0c3af: out <= 12'hb27;
      20'h0c3b0: out <= 12'hee9;
      20'h0c3b1: out <= 12'hf87;
      20'h0c3b2: out <= 12'hee9;
      20'h0c3b3: out <= 12'hee9;
      20'h0c3b4: out <= 12'hee9;
      20'h0c3b5: out <= 12'hb27;
      20'h0c3b6: out <= 12'hf87;
      20'h0c3b7: out <= 12'hb27;
      20'h0c3b8: out <= 12'hee9;
      20'h0c3b9: out <= 12'hf87;
      20'h0c3ba: out <= 12'hee9;
      20'h0c3bb: out <= 12'hee9;
      20'h0c3bc: out <= 12'hee9;
      20'h0c3bd: out <= 12'hb27;
      20'h0c3be: out <= 12'hf87;
      20'h0c3bf: out <= 12'hb27;
      20'h0c3c0: out <= 12'hee9;
      20'h0c3c1: out <= 12'hf87;
      20'h0c3c2: out <= 12'hee9;
      20'h0c3c3: out <= 12'hee9;
      20'h0c3c4: out <= 12'hee9;
      20'h0c3c5: out <= 12'hb27;
      20'h0c3c6: out <= 12'hf87;
      20'h0c3c7: out <= 12'hb27;
      20'h0c3c8: out <= 12'h088;
      20'h0c3c9: out <= 12'h088;
      20'h0c3ca: out <= 12'h088;
      20'h0c3cb: out <= 12'h088;
      20'h0c3cc: out <= 12'h088;
      20'h0c3cd: out <= 12'h088;
      20'h0c3ce: out <= 12'h088;
      20'h0c3cf: out <= 12'h088;
      20'h0c3d0: out <= 12'h088;
      20'h0c3d1: out <= 12'h088;
      20'h0c3d2: out <= 12'h088;
      20'h0c3d3: out <= 12'h088;
      20'h0c3d4: out <= 12'h088;
      20'h0c3d5: out <= 12'h088;
      20'h0c3d6: out <= 12'h088;
      20'h0c3d7: out <= 12'h088;
      20'h0c3d8: out <= 12'h088;
      20'h0c3d9: out <= 12'h088;
      20'h0c3da: out <= 12'h088;
      20'h0c3db: out <= 12'h088;
      20'h0c3dc: out <= 12'h088;
      20'h0c3dd: out <= 12'h088;
      20'h0c3de: out <= 12'h088;
      20'h0c3df: out <= 12'h088;
      20'h0c3e0: out <= 12'h088;
      20'h0c3e1: out <= 12'h088;
      20'h0c3e2: out <= 12'h088;
      20'h0c3e3: out <= 12'h088;
      20'h0c3e4: out <= 12'h088;
      20'h0c3e5: out <= 12'h088;
      20'h0c3e6: out <= 12'h088;
      20'h0c3e7: out <= 12'h088;
      20'h0c3e8: out <= 12'h088;
      20'h0c3e9: out <= 12'h088;
      20'h0c3ea: out <= 12'h088;
      20'h0c3eb: out <= 12'h088;
      20'h0c3ec: out <= 12'h088;
      20'h0c3ed: out <= 12'h088;
      20'h0c3ee: out <= 12'h088;
      20'h0c3ef: out <= 12'h088;
      20'h0c3f0: out <= 12'h088;
      20'h0c3f1: out <= 12'h088;
      20'h0c3f2: out <= 12'h088;
      20'h0c3f3: out <= 12'h088;
      20'h0c3f4: out <= 12'h088;
      20'h0c3f5: out <= 12'h088;
      20'h0c3f6: out <= 12'h088;
      20'h0c3f7: out <= 12'h088;
      20'h0c3f8: out <= 12'h088;
      20'h0c3f9: out <= 12'h088;
      20'h0c3fa: out <= 12'h088;
      20'h0c3fb: out <= 12'h088;
      20'h0c3fc: out <= 12'h088;
      20'h0c3fd: out <= 12'h088;
      20'h0c3fe: out <= 12'h088;
      20'h0c3ff: out <= 12'h088;
      20'h0c400: out <= 12'h088;
      20'h0c401: out <= 12'h088;
      20'h0c402: out <= 12'h088;
      20'h0c403: out <= 12'h088;
      20'h0c404: out <= 12'h088;
      20'h0c405: out <= 12'h088;
      20'h0c406: out <= 12'h088;
      20'h0c407: out <= 12'h088;
      20'h0c408: out <= 12'h088;
      20'h0c409: out <= 12'h088;
      20'h0c40a: out <= 12'h088;
      20'h0c40b: out <= 12'h088;
      20'h0c40c: out <= 12'h088;
      20'h0c40d: out <= 12'h088;
      20'h0c40e: out <= 12'h088;
      20'h0c40f: out <= 12'h088;
      20'h0c410: out <= 12'h088;
      20'h0c411: out <= 12'h088;
      20'h0c412: out <= 12'h088;
      20'h0c413: out <= 12'h088;
      20'h0c414: out <= 12'h088;
      20'h0c415: out <= 12'h088;
      20'h0c416: out <= 12'h088;
      20'h0c417: out <= 12'h088;
      20'h0c418: out <= 12'h088;
      20'h0c419: out <= 12'h088;
      20'h0c41a: out <= 12'h088;
      20'h0c41b: out <= 12'h088;
      20'h0c41c: out <= 12'h088;
      20'h0c41d: out <= 12'h088;
      20'h0c41e: out <= 12'h088;
      20'h0c41f: out <= 12'h088;
      20'h0c420: out <= 12'h088;
      20'h0c421: out <= 12'h088;
      20'h0c422: out <= 12'h088;
      20'h0c423: out <= 12'h088;
      20'h0c424: out <= 12'h088;
      20'h0c425: out <= 12'h088;
      20'h0c426: out <= 12'h088;
      20'h0c427: out <= 12'h088;
      20'h0c428: out <= 12'h088;
      20'h0c429: out <= 12'h088;
      20'h0c42a: out <= 12'h088;
      20'h0c42b: out <= 12'h088;
      20'h0c42c: out <= 12'h088;
      20'h0c42d: out <= 12'h088;
      20'h0c42e: out <= 12'h088;
      20'h0c42f: out <= 12'h088;
      20'h0c430: out <= 12'h088;
      20'h0c431: out <= 12'h222;
      20'h0c432: out <= 12'h222;
      20'h0c433: out <= 12'h222;
      20'h0c434: out <= 12'h222;
      20'h0c435: out <= 12'h222;
      20'h0c436: out <= 12'h222;
      20'h0c437: out <= 12'h222;
      20'h0c438: out <= 12'h660;
      20'h0c439: out <= 12'hbb0;
      20'h0c43a: out <= 12'hee9;
      20'h0c43b: out <= 12'hee9;
      20'h0c43c: out <= 12'hee9;
      20'h0c43d: out <= 12'hee9;
      20'h0c43e: out <= 12'hee9;
      20'h0c43f: out <= 12'hbb0;
      20'h0c440: out <= 12'h660;
      20'h0c441: out <= 12'h222;
      20'h0c442: out <= 12'h222;
      20'h0c443: out <= 12'h222;
      20'h0c444: out <= 12'h222;
      20'h0c445: out <= 12'h222;
      20'h0c446: out <= 12'h222;
      20'h0c447: out <= 12'h222;
      20'h0c448: out <= 12'h603;
      20'h0c449: out <= 12'h603;
      20'h0c44a: out <= 12'h603;
      20'h0c44b: out <= 12'h603;
      20'h0c44c: out <= 12'hf87;
      20'h0c44d: out <= 12'hf87;
      20'h0c44e: out <= 12'h000;
      20'h0c44f: out <= 12'h000;
      20'h0c450: out <= 12'h000;
      20'h0c451: out <= 12'hf87;
      20'h0c452: out <= 12'hf87;
      20'h0c453: out <= 12'h000;
      20'h0c454: out <= 12'h000;
      20'h0c455: out <= 12'h000;
      20'h0c456: out <= 12'h000;
      20'h0c457: out <= 12'hf87;
      20'h0c458: out <= 12'hf87;
      20'h0c459: out <= 12'h000;
      20'h0c45a: out <= 12'h000;
      20'h0c45b: out <= 12'h000;
      20'h0c45c: out <= 12'hf87;
      20'h0c45d: out <= 12'hf87;
      20'h0c45e: out <= 12'hf87;
      20'h0c45f: out <= 12'h000;
      20'h0c460: out <= 12'h000;
      20'h0c461: out <= 12'h000;
      20'h0c462: out <= 12'h000;
      20'h0c463: out <= 12'h000;
      20'h0c464: out <= 12'hf87;
      20'h0c465: out <= 12'hf87;
      20'h0c466: out <= 12'h000;
      20'h0c467: out <= 12'h000;
      20'h0c468: out <= 12'h000;
      20'h0c469: out <= 12'hf87;
      20'h0c46a: out <= 12'hf87;
      20'h0c46b: out <= 12'h000;
      20'h0c46c: out <= 12'hf87;
      20'h0c46d: out <= 12'hf87;
      20'h0c46e: out <= 12'hf87;
      20'h0c46f: out <= 12'hf87;
      20'h0c470: out <= 12'hf87;
      20'h0c471: out <= 12'hf87;
      20'h0c472: out <= 12'hf87;
      20'h0c473: out <= 12'h000;
      20'h0c474: out <= 12'hf87;
      20'h0c475: out <= 12'hf87;
      20'h0c476: out <= 12'h000;
      20'h0c477: out <= 12'h000;
      20'h0c478: out <= 12'h000;
      20'h0c479: out <= 12'hf87;
      20'h0c47a: out <= 12'hf87;
      20'h0c47b: out <= 12'h000;
      20'h0c47c: out <= 12'hf87;
      20'h0c47d: out <= 12'hf87;
      20'h0c47e: out <= 12'h000;
      20'h0c47f: out <= 12'h000;
      20'h0c480: out <= 12'h000;
      20'h0c481: out <= 12'hf87;
      20'h0c482: out <= 12'hf87;
      20'h0c483: out <= 12'h000;
      20'h0c484: out <= 12'h000;
      20'h0c485: out <= 12'h000;
      20'h0c486: out <= 12'hf87;
      20'h0c487: out <= 12'hf87;
      20'h0c488: out <= 12'h000;
      20'h0c489: out <= 12'h000;
      20'h0c48a: out <= 12'h000;
      20'h0c48b: out <= 12'h000;
      20'h0c48c: out <= 12'hf87;
      20'h0c48d: out <= 12'hf87;
      20'h0c48e: out <= 12'h000;
      20'h0c48f: out <= 12'h000;
      20'h0c490: out <= 12'h000;
      20'h0c491: out <= 12'hf87;
      20'h0c492: out <= 12'hf87;
      20'h0c493: out <= 12'h000;
      20'h0c494: out <= 12'h000;
      20'h0c495: out <= 12'h000;
      20'h0c496: out <= 12'h000;
      20'h0c497: out <= 12'hf87;
      20'h0c498: out <= 12'hf87;
      20'h0c499: out <= 12'hf87;
      20'h0c49a: out <= 12'h000;
      20'h0c49b: out <= 12'h000;
      20'h0c49c: out <= 12'h603;
      20'h0c49d: out <= 12'h603;
      20'h0c49e: out <= 12'h603;
      20'h0c49f: out <= 12'h603;
      20'h0c4a0: out <= 12'hee9;
      20'h0c4a1: out <= 12'hf87;
      20'h0c4a2: out <= 12'hee9;
      20'h0c4a3: out <= 12'hf87;
      20'h0c4a4: out <= 12'hf87;
      20'h0c4a5: out <= 12'hb27;
      20'h0c4a6: out <= 12'hf87;
      20'h0c4a7: out <= 12'hb27;
      20'h0c4a8: out <= 12'hee9;
      20'h0c4a9: out <= 12'hf87;
      20'h0c4aa: out <= 12'hee9;
      20'h0c4ab: out <= 12'hf87;
      20'h0c4ac: out <= 12'hf87;
      20'h0c4ad: out <= 12'hb27;
      20'h0c4ae: out <= 12'hf87;
      20'h0c4af: out <= 12'hb27;
      20'h0c4b0: out <= 12'hee9;
      20'h0c4b1: out <= 12'hf87;
      20'h0c4b2: out <= 12'hee9;
      20'h0c4b3: out <= 12'hf87;
      20'h0c4b4: out <= 12'hf87;
      20'h0c4b5: out <= 12'hb27;
      20'h0c4b6: out <= 12'hf87;
      20'h0c4b7: out <= 12'hb27;
      20'h0c4b8: out <= 12'hee9;
      20'h0c4b9: out <= 12'hf87;
      20'h0c4ba: out <= 12'hee9;
      20'h0c4bb: out <= 12'hf87;
      20'h0c4bc: out <= 12'hf87;
      20'h0c4bd: out <= 12'hb27;
      20'h0c4be: out <= 12'hf87;
      20'h0c4bf: out <= 12'hb27;
      20'h0c4c0: out <= 12'hee9;
      20'h0c4c1: out <= 12'hf87;
      20'h0c4c2: out <= 12'hee9;
      20'h0c4c3: out <= 12'hf87;
      20'h0c4c4: out <= 12'hf87;
      20'h0c4c5: out <= 12'hb27;
      20'h0c4c6: out <= 12'hf87;
      20'h0c4c7: out <= 12'hb27;
      20'h0c4c8: out <= 12'hee9;
      20'h0c4c9: out <= 12'hf87;
      20'h0c4ca: out <= 12'hee9;
      20'h0c4cb: out <= 12'hf87;
      20'h0c4cc: out <= 12'hf87;
      20'h0c4cd: out <= 12'hb27;
      20'h0c4ce: out <= 12'hf87;
      20'h0c4cf: out <= 12'hb27;
      20'h0c4d0: out <= 12'hee9;
      20'h0c4d1: out <= 12'hf87;
      20'h0c4d2: out <= 12'hee9;
      20'h0c4d3: out <= 12'hf87;
      20'h0c4d4: out <= 12'hf87;
      20'h0c4d5: out <= 12'hb27;
      20'h0c4d6: out <= 12'hf87;
      20'h0c4d7: out <= 12'hb27;
      20'h0c4d8: out <= 12'hee9;
      20'h0c4d9: out <= 12'hf87;
      20'h0c4da: out <= 12'hee9;
      20'h0c4db: out <= 12'hf87;
      20'h0c4dc: out <= 12'hf87;
      20'h0c4dd: out <= 12'hb27;
      20'h0c4de: out <= 12'hf87;
      20'h0c4df: out <= 12'hb27;
      20'h0c4e0: out <= 12'h088;
      20'h0c4e1: out <= 12'h088;
      20'h0c4e2: out <= 12'h088;
      20'h0c4e3: out <= 12'h088;
      20'h0c4e4: out <= 12'h088;
      20'h0c4e5: out <= 12'h088;
      20'h0c4e6: out <= 12'h088;
      20'h0c4e7: out <= 12'h088;
      20'h0c4e8: out <= 12'h088;
      20'h0c4e9: out <= 12'h088;
      20'h0c4ea: out <= 12'h088;
      20'h0c4eb: out <= 12'h088;
      20'h0c4ec: out <= 12'h088;
      20'h0c4ed: out <= 12'h088;
      20'h0c4ee: out <= 12'h088;
      20'h0c4ef: out <= 12'h088;
      20'h0c4f0: out <= 12'h088;
      20'h0c4f1: out <= 12'h088;
      20'h0c4f2: out <= 12'h088;
      20'h0c4f3: out <= 12'h088;
      20'h0c4f4: out <= 12'h088;
      20'h0c4f5: out <= 12'h088;
      20'h0c4f6: out <= 12'h088;
      20'h0c4f7: out <= 12'h088;
      20'h0c4f8: out <= 12'h088;
      20'h0c4f9: out <= 12'h088;
      20'h0c4fa: out <= 12'h088;
      20'h0c4fb: out <= 12'h088;
      20'h0c4fc: out <= 12'h088;
      20'h0c4fd: out <= 12'h088;
      20'h0c4fe: out <= 12'h088;
      20'h0c4ff: out <= 12'h088;
      20'h0c500: out <= 12'h088;
      20'h0c501: out <= 12'h088;
      20'h0c502: out <= 12'h088;
      20'h0c503: out <= 12'h088;
      20'h0c504: out <= 12'h088;
      20'h0c505: out <= 12'h088;
      20'h0c506: out <= 12'h088;
      20'h0c507: out <= 12'h088;
      20'h0c508: out <= 12'h088;
      20'h0c509: out <= 12'h088;
      20'h0c50a: out <= 12'h088;
      20'h0c50b: out <= 12'h088;
      20'h0c50c: out <= 12'h088;
      20'h0c50d: out <= 12'h088;
      20'h0c50e: out <= 12'h088;
      20'h0c50f: out <= 12'h088;
      20'h0c510: out <= 12'h088;
      20'h0c511: out <= 12'h088;
      20'h0c512: out <= 12'h088;
      20'h0c513: out <= 12'h088;
      20'h0c514: out <= 12'h088;
      20'h0c515: out <= 12'h088;
      20'h0c516: out <= 12'h088;
      20'h0c517: out <= 12'h088;
      20'h0c518: out <= 12'h088;
      20'h0c519: out <= 12'h088;
      20'h0c51a: out <= 12'h088;
      20'h0c51b: out <= 12'h088;
      20'h0c51c: out <= 12'h088;
      20'h0c51d: out <= 12'h088;
      20'h0c51e: out <= 12'h088;
      20'h0c51f: out <= 12'h088;
      20'h0c520: out <= 12'h088;
      20'h0c521: out <= 12'h088;
      20'h0c522: out <= 12'h088;
      20'h0c523: out <= 12'h088;
      20'h0c524: out <= 12'h088;
      20'h0c525: out <= 12'h088;
      20'h0c526: out <= 12'h088;
      20'h0c527: out <= 12'h088;
      20'h0c528: out <= 12'h088;
      20'h0c529: out <= 12'h088;
      20'h0c52a: out <= 12'h088;
      20'h0c52b: out <= 12'h088;
      20'h0c52c: out <= 12'h088;
      20'h0c52d: out <= 12'h088;
      20'h0c52e: out <= 12'h088;
      20'h0c52f: out <= 12'h088;
      20'h0c530: out <= 12'h088;
      20'h0c531: out <= 12'h088;
      20'h0c532: out <= 12'h088;
      20'h0c533: out <= 12'h088;
      20'h0c534: out <= 12'h088;
      20'h0c535: out <= 12'h088;
      20'h0c536: out <= 12'h088;
      20'h0c537: out <= 12'h088;
      20'h0c538: out <= 12'h088;
      20'h0c539: out <= 12'h088;
      20'h0c53a: out <= 12'h088;
      20'h0c53b: out <= 12'h088;
      20'h0c53c: out <= 12'h088;
      20'h0c53d: out <= 12'h088;
      20'h0c53e: out <= 12'h088;
      20'h0c53f: out <= 12'h088;
      20'h0c540: out <= 12'h088;
      20'h0c541: out <= 12'h088;
      20'h0c542: out <= 12'h088;
      20'h0c543: out <= 12'h088;
      20'h0c544: out <= 12'h088;
      20'h0c545: out <= 12'h088;
      20'h0c546: out <= 12'h088;
      20'h0c547: out <= 12'h088;
      20'h0c548: out <= 12'h088;
      20'h0c549: out <= 12'h222;
      20'h0c54a: out <= 12'h222;
      20'h0c54b: out <= 12'h222;
      20'h0c54c: out <= 12'h222;
      20'h0c54d: out <= 12'h222;
      20'h0c54e: out <= 12'h222;
      20'h0c54f: out <= 12'h222;
      20'h0c550: out <= 12'h222;
      20'h0c551: out <= 12'h660;
      20'h0c552: out <= 12'hbb0;
      20'h0c553: out <= 12'hee9;
      20'h0c554: out <= 12'hee9;
      20'h0c555: out <= 12'hee9;
      20'h0c556: out <= 12'hbb0;
      20'h0c557: out <= 12'h660;
      20'h0c558: out <= 12'h222;
      20'h0c559: out <= 12'h222;
      20'h0c55a: out <= 12'h222;
      20'h0c55b: out <= 12'h222;
      20'h0c55c: out <= 12'h222;
      20'h0c55d: out <= 12'h222;
      20'h0c55e: out <= 12'h222;
      20'h0c55f: out <= 12'h222;
      20'h0c560: out <= 12'h603;
      20'h0c561: out <= 12'h603;
      20'h0c562: out <= 12'h603;
      20'h0c563: out <= 12'h603;
      20'h0c564: out <= 12'hb27;
      20'h0c565: out <= 12'hb27;
      20'h0c566: out <= 12'hb27;
      20'h0c567: out <= 12'hb27;
      20'h0c568: out <= 12'hb27;
      20'h0c569: out <= 12'hb27;
      20'h0c56a: out <= 12'hb27;
      20'h0c56b: out <= 12'h000;
      20'h0c56c: out <= 12'h000;
      20'h0c56d: out <= 12'h000;
      20'h0c56e: out <= 12'h000;
      20'h0c56f: out <= 12'hb27;
      20'h0c570: out <= 12'hb27;
      20'h0c571: out <= 12'h000;
      20'h0c572: out <= 12'h000;
      20'h0c573: out <= 12'h000;
      20'h0c574: out <= 12'hb27;
      20'h0c575: out <= 12'hb27;
      20'h0c576: out <= 12'hb27;
      20'h0c577: out <= 12'hb27;
      20'h0c578: out <= 12'hb27;
      20'h0c579: out <= 12'hb27;
      20'h0c57a: out <= 12'hb27;
      20'h0c57b: out <= 12'h000;
      20'h0c57c: out <= 12'hb27;
      20'h0c57d: out <= 12'hb27;
      20'h0c57e: out <= 12'hb27;
      20'h0c57f: out <= 12'hb27;
      20'h0c580: out <= 12'hb27;
      20'h0c581: out <= 12'hb27;
      20'h0c582: out <= 12'hb27;
      20'h0c583: out <= 12'h000;
      20'h0c584: out <= 12'h000;
      20'h0c585: out <= 12'h000;
      20'h0c586: out <= 12'h000;
      20'h0c587: out <= 12'h000;
      20'h0c588: out <= 12'hb27;
      20'h0c589: out <= 12'hb27;
      20'h0c58a: out <= 12'h000;
      20'h0c58b: out <= 12'h000;
      20'h0c58c: out <= 12'hb27;
      20'h0c58d: out <= 12'hb27;
      20'h0c58e: out <= 12'hb27;
      20'h0c58f: out <= 12'hb27;
      20'h0c590: out <= 12'hb27;
      20'h0c591: out <= 12'hb27;
      20'h0c592: out <= 12'hb27;
      20'h0c593: out <= 12'h000;
      20'h0c594: out <= 12'hb27;
      20'h0c595: out <= 12'hb27;
      20'h0c596: out <= 12'hb27;
      20'h0c597: out <= 12'hb27;
      20'h0c598: out <= 12'hb27;
      20'h0c599: out <= 12'hb27;
      20'h0c59a: out <= 12'hb27;
      20'h0c59b: out <= 12'h000;
      20'h0c59c: out <= 12'h000;
      20'h0c59d: out <= 12'h000;
      20'h0c59e: out <= 12'hb27;
      20'h0c59f: out <= 12'hb27;
      20'h0c5a0: out <= 12'h000;
      20'h0c5a1: out <= 12'h000;
      20'h0c5a2: out <= 12'h000;
      20'h0c5a3: out <= 12'h000;
      20'h0c5a4: out <= 12'hb27;
      20'h0c5a5: out <= 12'hb27;
      20'h0c5a6: out <= 12'hb27;
      20'h0c5a7: out <= 12'hb27;
      20'h0c5a8: out <= 12'hb27;
      20'h0c5a9: out <= 12'hb27;
      20'h0c5aa: out <= 12'hb27;
      20'h0c5ab: out <= 12'h000;
      20'h0c5ac: out <= 12'h000;
      20'h0c5ad: out <= 12'hb27;
      20'h0c5ae: out <= 12'hb27;
      20'h0c5af: out <= 12'hb27;
      20'h0c5b0: out <= 12'hb27;
      20'h0c5b1: out <= 12'h000;
      20'h0c5b2: out <= 12'h000;
      20'h0c5b3: out <= 12'h000;
      20'h0c5b4: out <= 12'h603;
      20'h0c5b5: out <= 12'h603;
      20'h0c5b6: out <= 12'h603;
      20'h0c5b7: out <= 12'h603;
      20'h0c5b8: out <= 12'hee9;
      20'h0c5b9: out <= 12'hf87;
      20'h0c5ba: out <= 12'hee9;
      20'h0c5bb: out <= 12'hf87;
      20'h0c5bc: out <= 12'hf87;
      20'h0c5bd: out <= 12'hb27;
      20'h0c5be: out <= 12'hf87;
      20'h0c5bf: out <= 12'hb27;
      20'h0c5c0: out <= 12'hee9;
      20'h0c5c1: out <= 12'hf87;
      20'h0c5c2: out <= 12'hee9;
      20'h0c5c3: out <= 12'hf87;
      20'h0c5c4: out <= 12'hf87;
      20'h0c5c5: out <= 12'hb27;
      20'h0c5c6: out <= 12'hf87;
      20'h0c5c7: out <= 12'hb27;
      20'h0c5c8: out <= 12'hee9;
      20'h0c5c9: out <= 12'hf87;
      20'h0c5ca: out <= 12'hee9;
      20'h0c5cb: out <= 12'hf87;
      20'h0c5cc: out <= 12'hf87;
      20'h0c5cd: out <= 12'hb27;
      20'h0c5ce: out <= 12'hf87;
      20'h0c5cf: out <= 12'hb27;
      20'h0c5d0: out <= 12'hee9;
      20'h0c5d1: out <= 12'hf87;
      20'h0c5d2: out <= 12'hee9;
      20'h0c5d3: out <= 12'hf87;
      20'h0c5d4: out <= 12'hf87;
      20'h0c5d5: out <= 12'hb27;
      20'h0c5d6: out <= 12'hf87;
      20'h0c5d7: out <= 12'hb27;
      20'h0c5d8: out <= 12'hee9;
      20'h0c5d9: out <= 12'hf87;
      20'h0c5da: out <= 12'hee9;
      20'h0c5db: out <= 12'hf87;
      20'h0c5dc: out <= 12'hf87;
      20'h0c5dd: out <= 12'hb27;
      20'h0c5de: out <= 12'hf87;
      20'h0c5df: out <= 12'hb27;
      20'h0c5e0: out <= 12'hee9;
      20'h0c5e1: out <= 12'hf87;
      20'h0c5e2: out <= 12'hee9;
      20'h0c5e3: out <= 12'hf87;
      20'h0c5e4: out <= 12'hf87;
      20'h0c5e5: out <= 12'hb27;
      20'h0c5e6: out <= 12'hf87;
      20'h0c5e7: out <= 12'hb27;
      20'h0c5e8: out <= 12'hee9;
      20'h0c5e9: out <= 12'hf87;
      20'h0c5ea: out <= 12'hee9;
      20'h0c5eb: out <= 12'hf87;
      20'h0c5ec: out <= 12'hf87;
      20'h0c5ed: out <= 12'hb27;
      20'h0c5ee: out <= 12'hf87;
      20'h0c5ef: out <= 12'hb27;
      20'h0c5f0: out <= 12'hee9;
      20'h0c5f1: out <= 12'hf87;
      20'h0c5f2: out <= 12'hee9;
      20'h0c5f3: out <= 12'hf87;
      20'h0c5f4: out <= 12'hf87;
      20'h0c5f5: out <= 12'hb27;
      20'h0c5f6: out <= 12'hf87;
      20'h0c5f7: out <= 12'hb27;
      20'h0c5f8: out <= 12'h088;
      20'h0c5f9: out <= 12'h088;
      20'h0c5fa: out <= 12'h088;
      20'h0c5fb: out <= 12'h088;
      20'h0c5fc: out <= 12'h088;
      20'h0c5fd: out <= 12'h088;
      20'h0c5fe: out <= 12'h088;
      20'h0c5ff: out <= 12'h088;
      20'h0c600: out <= 12'h088;
      20'h0c601: out <= 12'h088;
      20'h0c602: out <= 12'h088;
      20'h0c603: out <= 12'h088;
      20'h0c604: out <= 12'h088;
      20'h0c605: out <= 12'h088;
      20'h0c606: out <= 12'h088;
      20'h0c607: out <= 12'h088;
      20'h0c608: out <= 12'h088;
      20'h0c609: out <= 12'h088;
      20'h0c60a: out <= 12'h088;
      20'h0c60b: out <= 12'h088;
      20'h0c60c: out <= 12'h088;
      20'h0c60d: out <= 12'h088;
      20'h0c60e: out <= 12'h088;
      20'h0c60f: out <= 12'h088;
      20'h0c610: out <= 12'h088;
      20'h0c611: out <= 12'h088;
      20'h0c612: out <= 12'h088;
      20'h0c613: out <= 12'h088;
      20'h0c614: out <= 12'h088;
      20'h0c615: out <= 12'h088;
      20'h0c616: out <= 12'h088;
      20'h0c617: out <= 12'h088;
      20'h0c618: out <= 12'h088;
      20'h0c619: out <= 12'h088;
      20'h0c61a: out <= 12'h088;
      20'h0c61b: out <= 12'h088;
      20'h0c61c: out <= 12'h088;
      20'h0c61d: out <= 12'h088;
      20'h0c61e: out <= 12'h088;
      20'h0c61f: out <= 12'h088;
      20'h0c620: out <= 12'h088;
      20'h0c621: out <= 12'h088;
      20'h0c622: out <= 12'h088;
      20'h0c623: out <= 12'h088;
      20'h0c624: out <= 12'h088;
      20'h0c625: out <= 12'h088;
      20'h0c626: out <= 12'h088;
      20'h0c627: out <= 12'h088;
      20'h0c628: out <= 12'h088;
      20'h0c629: out <= 12'h088;
      20'h0c62a: out <= 12'h088;
      20'h0c62b: out <= 12'h088;
      20'h0c62c: out <= 12'h088;
      20'h0c62d: out <= 12'h088;
      20'h0c62e: out <= 12'h088;
      20'h0c62f: out <= 12'h088;
      20'h0c630: out <= 12'h088;
      20'h0c631: out <= 12'h088;
      20'h0c632: out <= 12'h088;
      20'h0c633: out <= 12'h088;
      20'h0c634: out <= 12'h088;
      20'h0c635: out <= 12'h088;
      20'h0c636: out <= 12'h088;
      20'h0c637: out <= 12'h088;
      20'h0c638: out <= 12'h088;
      20'h0c639: out <= 12'h088;
      20'h0c63a: out <= 12'h088;
      20'h0c63b: out <= 12'h088;
      20'h0c63c: out <= 12'h088;
      20'h0c63d: out <= 12'h088;
      20'h0c63e: out <= 12'h088;
      20'h0c63f: out <= 12'h088;
      20'h0c640: out <= 12'h088;
      20'h0c641: out <= 12'h088;
      20'h0c642: out <= 12'h088;
      20'h0c643: out <= 12'h088;
      20'h0c644: out <= 12'h088;
      20'h0c645: out <= 12'h088;
      20'h0c646: out <= 12'h088;
      20'h0c647: out <= 12'h088;
      20'h0c648: out <= 12'h088;
      20'h0c649: out <= 12'h088;
      20'h0c64a: out <= 12'h088;
      20'h0c64b: out <= 12'h088;
      20'h0c64c: out <= 12'h088;
      20'h0c64d: out <= 12'h088;
      20'h0c64e: out <= 12'h088;
      20'h0c64f: out <= 12'h088;
      20'h0c650: out <= 12'h088;
      20'h0c651: out <= 12'h088;
      20'h0c652: out <= 12'h088;
      20'h0c653: out <= 12'h088;
      20'h0c654: out <= 12'h088;
      20'h0c655: out <= 12'h088;
      20'h0c656: out <= 12'h088;
      20'h0c657: out <= 12'h088;
      20'h0c658: out <= 12'h088;
      20'h0c659: out <= 12'h088;
      20'h0c65a: out <= 12'h088;
      20'h0c65b: out <= 12'h088;
      20'h0c65c: out <= 12'h088;
      20'h0c65d: out <= 12'h088;
      20'h0c65e: out <= 12'h088;
      20'h0c65f: out <= 12'h088;
      20'h0c660: out <= 12'h088;
      20'h0c661: out <= 12'h222;
      20'h0c662: out <= 12'h222;
      20'h0c663: out <= 12'h222;
      20'h0c664: out <= 12'h222;
      20'h0c665: out <= 12'h222;
      20'h0c666: out <= 12'h222;
      20'h0c667: out <= 12'h222;
      20'h0c668: out <= 12'h222;
      20'h0c669: out <= 12'h222;
      20'h0c66a: out <= 12'h660;
      20'h0c66b: out <= 12'hbb0;
      20'h0c66c: out <= 12'hee9;
      20'h0c66d: out <= 12'hbb0;
      20'h0c66e: out <= 12'h660;
      20'h0c66f: out <= 12'h222;
      20'h0c670: out <= 12'h222;
      20'h0c671: out <= 12'h222;
      20'h0c672: out <= 12'h222;
      20'h0c673: out <= 12'h222;
      20'h0c674: out <= 12'h222;
      20'h0c675: out <= 12'h222;
      20'h0c676: out <= 12'h222;
      20'h0c677: out <= 12'h222;
      20'h0c678: out <= 12'h603;
      20'h0c679: out <= 12'h603;
      20'h0c67a: out <= 12'h603;
      20'h0c67b: out <= 12'h603;
      20'h0c67c: out <= 12'h000;
      20'h0c67d: out <= 12'hb27;
      20'h0c67e: out <= 12'hb27;
      20'h0c67f: out <= 12'hb27;
      20'h0c680: out <= 12'hb27;
      20'h0c681: out <= 12'hb27;
      20'h0c682: out <= 12'h000;
      20'h0c683: out <= 12'h000;
      20'h0c684: out <= 12'h000;
      20'h0c685: out <= 12'h000;
      20'h0c686: out <= 12'h000;
      20'h0c687: out <= 12'hb27;
      20'h0c688: out <= 12'hb27;
      20'h0c689: out <= 12'h000;
      20'h0c68a: out <= 12'h000;
      20'h0c68b: out <= 12'h000;
      20'h0c68c: out <= 12'hb27;
      20'h0c68d: out <= 12'hb27;
      20'h0c68e: out <= 12'hb27;
      20'h0c68f: out <= 12'hb27;
      20'h0c690: out <= 12'hb27;
      20'h0c691: out <= 12'hb27;
      20'h0c692: out <= 12'hb27;
      20'h0c693: out <= 12'h000;
      20'h0c694: out <= 12'h000;
      20'h0c695: out <= 12'hb27;
      20'h0c696: out <= 12'hb27;
      20'h0c697: out <= 12'hb27;
      20'h0c698: out <= 12'hb27;
      20'h0c699: out <= 12'hb27;
      20'h0c69a: out <= 12'h000;
      20'h0c69b: out <= 12'h000;
      20'h0c69c: out <= 12'h000;
      20'h0c69d: out <= 12'h000;
      20'h0c69e: out <= 12'h000;
      20'h0c69f: out <= 12'h000;
      20'h0c6a0: out <= 12'hb27;
      20'h0c6a1: out <= 12'hb27;
      20'h0c6a2: out <= 12'h000;
      20'h0c6a3: out <= 12'h000;
      20'h0c6a4: out <= 12'h000;
      20'h0c6a5: out <= 12'hb27;
      20'h0c6a6: out <= 12'hb27;
      20'h0c6a7: out <= 12'hb27;
      20'h0c6a8: out <= 12'hb27;
      20'h0c6a9: out <= 12'hb27;
      20'h0c6aa: out <= 12'h000;
      20'h0c6ab: out <= 12'h000;
      20'h0c6ac: out <= 12'h000;
      20'h0c6ad: out <= 12'hb27;
      20'h0c6ae: out <= 12'hb27;
      20'h0c6af: out <= 12'hb27;
      20'h0c6b0: out <= 12'hb27;
      20'h0c6b1: out <= 12'hb27;
      20'h0c6b2: out <= 12'h000;
      20'h0c6b3: out <= 12'h000;
      20'h0c6b4: out <= 12'h000;
      20'h0c6b5: out <= 12'h000;
      20'h0c6b6: out <= 12'hb27;
      20'h0c6b7: out <= 12'hb27;
      20'h0c6b8: out <= 12'h000;
      20'h0c6b9: out <= 12'h000;
      20'h0c6ba: out <= 12'h000;
      20'h0c6bb: out <= 12'h000;
      20'h0c6bc: out <= 12'h000;
      20'h0c6bd: out <= 12'hb27;
      20'h0c6be: out <= 12'hb27;
      20'h0c6bf: out <= 12'hb27;
      20'h0c6c0: out <= 12'hb27;
      20'h0c6c1: out <= 12'hb27;
      20'h0c6c2: out <= 12'h000;
      20'h0c6c3: out <= 12'h000;
      20'h0c6c4: out <= 12'h000;
      20'h0c6c5: out <= 12'hb27;
      20'h0c6c6: out <= 12'hb27;
      20'h0c6c7: out <= 12'hb27;
      20'h0c6c8: out <= 12'h000;
      20'h0c6c9: out <= 12'h000;
      20'h0c6ca: out <= 12'h000;
      20'h0c6cb: out <= 12'h000;
      20'h0c6cc: out <= 12'h603;
      20'h0c6cd: out <= 12'h603;
      20'h0c6ce: out <= 12'h603;
      20'h0c6cf: out <= 12'h603;
      20'h0c6d0: out <= 12'hee9;
      20'h0c6d1: out <= 12'hf87;
      20'h0c6d2: out <= 12'hee9;
      20'h0c6d3: out <= 12'hb27;
      20'h0c6d4: out <= 12'hb27;
      20'h0c6d5: out <= 12'hb27;
      20'h0c6d6: out <= 12'hf87;
      20'h0c6d7: out <= 12'hb27;
      20'h0c6d8: out <= 12'hee9;
      20'h0c6d9: out <= 12'hf87;
      20'h0c6da: out <= 12'hee9;
      20'h0c6db: out <= 12'hb27;
      20'h0c6dc: out <= 12'hb27;
      20'h0c6dd: out <= 12'hb27;
      20'h0c6de: out <= 12'hf87;
      20'h0c6df: out <= 12'hb27;
      20'h0c6e0: out <= 12'hee9;
      20'h0c6e1: out <= 12'hf87;
      20'h0c6e2: out <= 12'hee9;
      20'h0c6e3: out <= 12'hb27;
      20'h0c6e4: out <= 12'hb27;
      20'h0c6e5: out <= 12'hb27;
      20'h0c6e6: out <= 12'hf87;
      20'h0c6e7: out <= 12'hb27;
      20'h0c6e8: out <= 12'hee9;
      20'h0c6e9: out <= 12'hf87;
      20'h0c6ea: out <= 12'hee9;
      20'h0c6eb: out <= 12'hb27;
      20'h0c6ec: out <= 12'hb27;
      20'h0c6ed: out <= 12'hb27;
      20'h0c6ee: out <= 12'hf87;
      20'h0c6ef: out <= 12'hb27;
      20'h0c6f0: out <= 12'hee9;
      20'h0c6f1: out <= 12'hf87;
      20'h0c6f2: out <= 12'hee9;
      20'h0c6f3: out <= 12'hb27;
      20'h0c6f4: out <= 12'hb27;
      20'h0c6f5: out <= 12'hb27;
      20'h0c6f6: out <= 12'hf87;
      20'h0c6f7: out <= 12'hb27;
      20'h0c6f8: out <= 12'hee9;
      20'h0c6f9: out <= 12'hf87;
      20'h0c6fa: out <= 12'hee9;
      20'h0c6fb: out <= 12'hb27;
      20'h0c6fc: out <= 12'hb27;
      20'h0c6fd: out <= 12'hb27;
      20'h0c6fe: out <= 12'hf87;
      20'h0c6ff: out <= 12'hb27;
      20'h0c700: out <= 12'hee9;
      20'h0c701: out <= 12'hf87;
      20'h0c702: out <= 12'hee9;
      20'h0c703: out <= 12'hb27;
      20'h0c704: out <= 12'hb27;
      20'h0c705: out <= 12'hb27;
      20'h0c706: out <= 12'hf87;
      20'h0c707: out <= 12'hb27;
      20'h0c708: out <= 12'hee9;
      20'h0c709: out <= 12'hf87;
      20'h0c70a: out <= 12'hee9;
      20'h0c70b: out <= 12'hb27;
      20'h0c70c: out <= 12'hb27;
      20'h0c70d: out <= 12'hb27;
      20'h0c70e: out <= 12'hf87;
      20'h0c70f: out <= 12'hb27;
      20'h0c710: out <= 12'h088;
      20'h0c711: out <= 12'h088;
      20'h0c712: out <= 12'h088;
      20'h0c713: out <= 12'h088;
      20'h0c714: out <= 12'h088;
      20'h0c715: out <= 12'h088;
      20'h0c716: out <= 12'h088;
      20'h0c717: out <= 12'h088;
      20'h0c718: out <= 12'h088;
      20'h0c719: out <= 12'h088;
      20'h0c71a: out <= 12'h088;
      20'h0c71b: out <= 12'h088;
      20'h0c71c: out <= 12'h088;
      20'h0c71d: out <= 12'h088;
      20'h0c71e: out <= 12'h088;
      20'h0c71f: out <= 12'h088;
      20'h0c720: out <= 12'h088;
      20'h0c721: out <= 12'h088;
      20'h0c722: out <= 12'h088;
      20'h0c723: out <= 12'h088;
      20'h0c724: out <= 12'h088;
      20'h0c725: out <= 12'h088;
      20'h0c726: out <= 12'h088;
      20'h0c727: out <= 12'h088;
      20'h0c728: out <= 12'h088;
      20'h0c729: out <= 12'h088;
      20'h0c72a: out <= 12'h088;
      20'h0c72b: out <= 12'h088;
      20'h0c72c: out <= 12'h088;
      20'h0c72d: out <= 12'h088;
      20'h0c72e: out <= 12'h088;
      20'h0c72f: out <= 12'h088;
      20'h0c730: out <= 12'h088;
      20'h0c731: out <= 12'h088;
      20'h0c732: out <= 12'h088;
      20'h0c733: out <= 12'h088;
      20'h0c734: out <= 12'h088;
      20'h0c735: out <= 12'h088;
      20'h0c736: out <= 12'h088;
      20'h0c737: out <= 12'h088;
      20'h0c738: out <= 12'h088;
      20'h0c739: out <= 12'h088;
      20'h0c73a: out <= 12'h088;
      20'h0c73b: out <= 12'h088;
      20'h0c73c: out <= 12'h088;
      20'h0c73d: out <= 12'h088;
      20'h0c73e: out <= 12'h088;
      20'h0c73f: out <= 12'h088;
      20'h0c740: out <= 12'h088;
      20'h0c741: out <= 12'h088;
      20'h0c742: out <= 12'h088;
      20'h0c743: out <= 12'h088;
      20'h0c744: out <= 12'h088;
      20'h0c745: out <= 12'h088;
      20'h0c746: out <= 12'h088;
      20'h0c747: out <= 12'h088;
      20'h0c748: out <= 12'h088;
      20'h0c749: out <= 12'h088;
      20'h0c74a: out <= 12'h088;
      20'h0c74b: out <= 12'h088;
      20'h0c74c: out <= 12'h088;
      20'h0c74d: out <= 12'h088;
      20'h0c74e: out <= 12'h088;
      20'h0c74f: out <= 12'h088;
      20'h0c750: out <= 12'h088;
      20'h0c751: out <= 12'h088;
      20'h0c752: out <= 12'h088;
      20'h0c753: out <= 12'h088;
      20'h0c754: out <= 12'h088;
      20'h0c755: out <= 12'h088;
      20'h0c756: out <= 12'h088;
      20'h0c757: out <= 12'h088;
      20'h0c758: out <= 12'h088;
      20'h0c759: out <= 12'h088;
      20'h0c75a: out <= 12'h088;
      20'h0c75b: out <= 12'h088;
      20'h0c75c: out <= 12'h088;
      20'h0c75d: out <= 12'h088;
      20'h0c75e: out <= 12'h088;
      20'h0c75f: out <= 12'h088;
      20'h0c760: out <= 12'h088;
      20'h0c761: out <= 12'h088;
      20'h0c762: out <= 12'h088;
      20'h0c763: out <= 12'h088;
      20'h0c764: out <= 12'h088;
      20'h0c765: out <= 12'h088;
      20'h0c766: out <= 12'h088;
      20'h0c767: out <= 12'h088;
      20'h0c768: out <= 12'h088;
      20'h0c769: out <= 12'h088;
      20'h0c76a: out <= 12'h088;
      20'h0c76b: out <= 12'h088;
      20'h0c76c: out <= 12'h088;
      20'h0c76d: out <= 12'h088;
      20'h0c76e: out <= 12'h088;
      20'h0c76f: out <= 12'h088;
      20'h0c770: out <= 12'h088;
      20'h0c771: out <= 12'h088;
      20'h0c772: out <= 12'h088;
      20'h0c773: out <= 12'h088;
      20'h0c774: out <= 12'h088;
      20'h0c775: out <= 12'h088;
      20'h0c776: out <= 12'h088;
      20'h0c777: out <= 12'h088;
      20'h0c778: out <= 12'h088;
      20'h0c779: out <= 12'h222;
      20'h0c77a: out <= 12'h222;
      20'h0c77b: out <= 12'h222;
      20'h0c77c: out <= 12'h222;
      20'h0c77d: out <= 12'h222;
      20'h0c77e: out <= 12'h222;
      20'h0c77f: out <= 12'h222;
      20'h0c780: out <= 12'h222;
      20'h0c781: out <= 12'h222;
      20'h0c782: out <= 12'h222;
      20'h0c783: out <= 12'h660;
      20'h0c784: out <= 12'hee9;
      20'h0c785: out <= 12'h660;
      20'h0c786: out <= 12'h222;
      20'h0c787: out <= 12'h222;
      20'h0c788: out <= 12'h222;
      20'h0c789: out <= 12'h222;
      20'h0c78a: out <= 12'h222;
      20'h0c78b: out <= 12'h222;
      20'h0c78c: out <= 12'h222;
      20'h0c78d: out <= 12'h222;
      20'h0c78e: out <= 12'h222;
      20'h0c78f: out <= 12'h222;
      20'h0c790: out <= 12'h603;
      20'h0c791: out <= 12'h603;
      20'h0c792: out <= 12'h603;
      20'h0c793: out <= 12'h603;
      20'h0c794: out <= 12'h000;
      20'h0c795: out <= 12'h000;
      20'h0c796: out <= 12'h000;
      20'h0c797: out <= 12'h000;
      20'h0c798: out <= 12'h000;
      20'h0c799: out <= 12'h000;
      20'h0c79a: out <= 12'h000;
      20'h0c79b: out <= 12'h000;
      20'h0c79c: out <= 12'h000;
      20'h0c79d: out <= 12'h000;
      20'h0c79e: out <= 12'h000;
      20'h0c79f: out <= 12'h000;
      20'h0c7a0: out <= 12'h000;
      20'h0c7a1: out <= 12'h000;
      20'h0c7a2: out <= 12'h000;
      20'h0c7a3: out <= 12'h000;
      20'h0c7a4: out <= 12'h000;
      20'h0c7a5: out <= 12'h000;
      20'h0c7a6: out <= 12'h000;
      20'h0c7a7: out <= 12'h000;
      20'h0c7a8: out <= 12'h000;
      20'h0c7a9: out <= 12'h000;
      20'h0c7aa: out <= 12'h000;
      20'h0c7ab: out <= 12'h000;
      20'h0c7ac: out <= 12'h000;
      20'h0c7ad: out <= 12'h000;
      20'h0c7ae: out <= 12'h000;
      20'h0c7af: out <= 12'h000;
      20'h0c7b0: out <= 12'h000;
      20'h0c7b1: out <= 12'h000;
      20'h0c7b2: out <= 12'h000;
      20'h0c7b3: out <= 12'h000;
      20'h0c7b4: out <= 12'h000;
      20'h0c7b5: out <= 12'h000;
      20'h0c7b6: out <= 12'h000;
      20'h0c7b7: out <= 12'h000;
      20'h0c7b8: out <= 12'h000;
      20'h0c7b9: out <= 12'h000;
      20'h0c7ba: out <= 12'h000;
      20'h0c7bb: out <= 12'h000;
      20'h0c7bc: out <= 12'h000;
      20'h0c7bd: out <= 12'h000;
      20'h0c7be: out <= 12'h000;
      20'h0c7bf: out <= 12'h000;
      20'h0c7c0: out <= 12'h000;
      20'h0c7c1: out <= 12'h000;
      20'h0c7c2: out <= 12'h000;
      20'h0c7c3: out <= 12'h000;
      20'h0c7c4: out <= 12'h000;
      20'h0c7c5: out <= 12'h000;
      20'h0c7c6: out <= 12'h000;
      20'h0c7c7: out <= 12'h000;
      20'h0c7c8: out <= 12'h000;
      20'h0c7c9: out <= 12'h000;
      20'h0c7ca: out <= 12'h000;
      20'h0c7cb: out <= 12'h000;
      20'h0c7cc: out <= 12'h000;
      20'h0c7cd: out <= 12'h000;
      20'h0c7ce: out <= 12'h000;
      20'h0c7cf: out <= 12'h000;
      20'h0c7d0: out <= 12'h000;
      20'h0c7d1: out <= 12'h000;
      20'h0c7d2: out <= 12'h000;
      20'h0c7d3: out <= 12'h000;
      20'h0c7d4: out <= 12'h000;
      20'h0c7d5: out <= 12'h000;
      20'h0c7d6: out <= 12'h000;
      20'h0c7d7: out <= 12'h000;
      20'h0c7d8: out <= 12'h000;
      20'h0c7d9: out <= 12'h000;
      20'h0c7da: out <= 12'h000;
      20'h0c7db: out <= 12'h000;
      20'h0c7dc: out <= 12'h000;
      20'h0c7dd: out <= 12'h000;
      20'h0c7de: out <= 12'h000;
      20'h0c7df: out <= 12'h000;
      20'h0c7e0: out <= 12'h000;
      20'h0c7e1: out <= 12'h000;
      20'h0c7e2: out <= 12'h000;
      20'h0c7e3: out <= 12'h000;
      20'h0c7e4: out <= 12'h603;
      20'h0c7e5: out <= 12'h603;
      20'h0c7e6: out <= 12'h603;
      20'h0c7e7: out <= 12'h603;
      20'h0c7e8: out <= 12'hee9;
      20'h0c7e9: out <= 12'hf87;
      20'h0c7ea: out <= 12'hf87;
      20'h0c7eb: out <= 12'hf87;
      20'h0c7ec: out <= 12'hf87;
      20'h0c7ed: out <= 12'hf87;
      20'h0c7ee: out <= 12'hf87;
      20'h0c7ef: out <= 12'hb27;
      20'h0c7f0: out <= 12'hee9;
      20'h0c7f1: out <= 12'hf87;
      20'h0c7f2: out <= 12'hf87;
      20'h0c7f3: out <= 12'hf87;
      20'h0c7f4: out <= 12'hf87;
      20'h0c7f5: out <= 12'hf87;
      20'h0c7f6: out <= 12'hf87;
      20'h0c7f7: out <= 12'hb27;
      20'h0c7f8: out <= 12'hee9;
      20'h0c7f9: out <= 12'hf87;
      20'h0c7fa: out <= 12'hf87;
      20'h0c7fb: out <= 12'hf87;
      20'h0c7fc: out <= 12'hf87;
      20'h0c7fd: out <= 12'hf87;
      20'h0c7fe: out <= 12'hf87;
      20'h0c7ff: out <= 12'hb27;
      20'h0c800: out <= 12'hee9;
      20'h0c801: out <= 12'hf87;
      20'h0c802: out <= 12'hf87;
      20'h0c803: out <= 12'hf87;
      20'h0c804: out <= 12'hf87;
      20'h0c805: out <= 12'hf87;
      20'h0c806: out <= 12'hf87;
      20'h0c807: out <= 12'hb27;
      20'h0c808: out <= 12'hee9;
      20'h0c809: out <= 12'hf87;
      20'h0c80a: out <= 12'hf87;
      20'h0c80b: out <= 12'hf87;
      20'h0c80c: out <= 12'hf87;
      20'h0c80d: out <= 12'hf87;
      20'h0c80e: out <= 12'hf87;
      20'h0c80f: out <= 12'hb27;
      20'h0c810: out <= 12'hee9;
      20'h0c811: out <= 12'hf87;
      20'h0c812: out <= 12'hf87;
      20'h0c813: out <= 12'hf87;
      20'h0c814: out <= 12'hf87;
      20'h0c815: out <= 12'hf87;
      20'h0c816: out <= 12'hf87;
      20'h0c817: out <= 12'hb27;
      20'h0c818: out <= 12'hee9;
      20'h0c819: out <= 12'hf87;
      20'h0c81a: out <= 12'hf87;
      20'h0c81b: out <= 12'hf87;
      20'h0c81c: out <= 12'hf87;
      20'h0c81d: out <= 12'hf87;
      20'h0c81e: out <= 12'hf87;
      20'h0c81f: out <= 12'hb27;
      20'h0c820: out <= 12'hee9;
      20'h0c821: out <= 12'hf87;
      20'h0c822: out <= 12'hf87;
      20'h0c823: out <= 12'hf87;
      20'h0c824: out <= 12'hf87;
      20'h0c825: out <= 12'hf87;
      20'h0c826: out <= 12'hf87;
      20'h0c827: out <= 12'hb27;
      20'h0c828: out <= 12'h088;
      20'h0c829: out <= 12'h088;
      20'h0c82a: out <= 12'h088;
      20'h0c82b: out <= 12'h088;
      20'h0c82c: out <= 12'h088;
      20'h0c82d: out <= 12'h088;
      20'h0c82e: out <= 12'h088;
      20'h0c82f: out <= 12'h088;
      20'h0c830: out <= 12'h088;
      20'h0c831: out <= 12'h088;
      20'h0c832: out <= 12'h088;
      20'h0c833: out <= 12'h088;
      20'h0c834: out <= 12'h088;
      20'h0c835: out <= 12'h088;
      20'h0c836: out <= 12'h088;
      20'h0c837: out <= 12'h088;
      20'h0c838: out <= 12'h088;
      20'h0c839: out <= 12'h088;
      20'h0c83a: out <= 12'h088;
      20'h0c83b: out <= 12'h088;
      20'h0c83c: out <= 12'h088;
      20'h0c83d: out <= 12'h088;
      20'h0c83e: out <= 12'h088;
      20'h0c83f: out <= 12'h088;
      20'h0c840: out <= 12'h088;
      20'h0c841: out <= 12'h088;
      20'h0c842: out <= 12'h088;
      20'h0c843: out <= 12'h088;
      20'h0c844: out <= 12'h088;
      20'h0c845: out <= 12'h088;
      20'h0c846: out <= 12'h088;
      20'h0c847: out <= 12'h088;
      20'h0c848: out <= 12'h088;
      20'h0c849: out <= 12'h088;
      20'h0c84a: out <= 12'h088;
      20'h0c84b: out <= 12'h088;
      20'h0c84c: out <= 12'h088;
      20'h0c84d: out <= 12'h088;
      20'h0c84e: out <= 12'h088;
      20'h0c84f: out <= 12'h088;
      20'h0c850: out <= 12'h088;
      20'h0c851: out <= 12'h088;
      20'h0c852: out <= 12'h088;
      20'h0c853: out <= 12'h088;
      20'h0c854: out <= 12'h088;
      20'h0c855: out <= 12'h088;
      20'h0c856: out <= 12'h088;
      20'h0c857: out <= 12'h088;
      20'h0c858: out <= 12'h088;
      20'h0c859: out <= 12'h088;
      20'h0c85a: out <= 12'h088;
      20'h0c85b: out <= 12'h088;
      20'h0c85c: out <= 12'h088;
      20'h0c85d: out <= 12'h088;
      20'h0c85e: out <= 12'h088;
      20'h0c85f: out <= 12'h088;
      20'h0c860: out <= 12'h088;
      20'h0c861: out <= 12'h088;
      20'h0c862: out <= 12'h088;
      20'h0c863: out <= 12'h088;
      20'h0c864: out <= 12'h088;
      20'h0c865: out <= 12'h088;
      20'h0c866: out <= 12'h088;
      20'h0c867: out <= 12'h088;
      20'h0c868: out <= 12'h088;
      20'h0c869: out <= 12'h088;
      20'h0c86a: out <= 12'h088;
      20'h0c86b: out <= 12'h088;
      20'h0c86c: out <= 12'h088;
      20'h0c86d: out <= 12'h088;
      20'h0c86e: out <= 12'h088;
      20'h0c86f: out <= 12'h088;
      20'h0c870: out <= 12'h088;
      20'h0c871: out <= 12'h088;
      20'h0c872: out <= 12'h088;
      20'h0c873: out <= 12'h088;
      20'h0c874: out <= 12'h088;
      20'h0c875: out <= 12'h088;
      20'h0c876: out <= 12'h088;
      20'h0c877: out <= 12'h088;
      20'h0c878: out <= 12'h088;
      20'h0c879: out <= 12'h088;
      20'h0c87a: out <= 12'h088;
      20'h0c87b: out <= 12'h088;
      20'h0c87c: out <= 12'h088;
      20'h0c87d: out <= 12'h088;
      20'h0c87e: out <= 12'h088;
      20'h0c87f: out <= 12'h088;
      20'h0c880: out <= 12'h088;
      20'h0c881: out <= 12'h088;
      20'h0c882: out <= 12'h088;
      20'h0c883: out <= 12'h088;
      20'h0c884: out <= 12'h088;
      20'h0c885: out <= 12'h088;
      20'h0c886: out <= 12'h088;
      20'h0c887: out <= 12'h088;
      20'h0c888: out <= 12'h088;
      20'h0c889: out <= 12'h088;
      20'h0c88a: out <= 12'h088;
      20'h0c88b: out <= 12'h088;
      20'h0c88c: out <= 12'h088;
      20'h0c88d: out <= 12'h088;
      20'h0c88e: out <= 12'h088;
      20'h0c88f: out <= 12'h088;
      20'h0c890: out <= 12'h088;
      20'h0c891: out <= 12'h222;
      20'h0c892: out <= 12'h222;
      20'h0c893: out <= 12'h222;
      20'h0c894: out <= 12'h222;
      20'h0c895: out <= 12'h222;
      20'h0c896: out <= 12'h222;
      20'h0c897: out <= 12'h222;
      20'h0c898: out <= 12'h222;
      20'h0c899: out <= 12'h222;
      20'h0c89a: out <= 12'h222;
      20'h0c89b: out <= 12'h222;
      20'h0c89c: out <= 12'hbb0;
      20'h0c89d: out <= 12'h222;
      20'h0c89e: out <= 12'h222;
      20'h0c89f: out <= 12'h222;
      20'h0c8a0: out <= 12'h222;
      20'h0c8a1: out <= 12'h222;
      20'h0c8a2: out <= 12'h222;
      20'h0c8a3: out <= 12'h222;
      20'h0c8a4: out <= 12'h222;
      20'h0c8a5: out <= 12'h222;
      20'h0c8a6: out <= 12'h222;
      20'h0c8a7: out <= 12'h222;
      20'h0c8a8: out <= 12'h603;
      20'h0c8a9: out <= 12'h603;
      20'h0c8aa: out <= 12'h603;
      20'h0c8ab: out <= 12'h603;
      20'h0c8ac: out <= 12'h000;
      20'h0c8ad: out <= 12'h000;
      20'h0c8ae: out <= 12'h000;
      20'h0c8af: out <= 12'h000;
      20'h0c8b0: out <= 12'h000;
      20'h0c8b1: out <= 12'h000;
      20'h0c8b2: out <= 12'h000;
      20'h0c8b3: out <= 12'h000;
      20'h0c8b4: out <= 12'h000;
      20'h0c8b5: out <= 12'h000;
      20'h0c8b6: out <= 12'h000;
      20'h0c8b7: out <= 12'h000;
      20'h0c8b8: out <= 12'h000;
      20'h0c8b9: out <= 12'h000;
      20'h0c8ba: out <= 12'h000;
      20'h0c8bb: out <= 12'h000;
      20'h0c8bc: out <= 12'h000;
      20'h0c8bd: out <= 12'h000;
      20'h0c8be: out <= 12'h000;
      20'h0c8bf: out <= 12'h000;
      20'h0c8c0: out <= 12'h000;
      20'h0c8c1: out <= 12'h000;
      20'h0c8c2: out <= 12'h000;
      20'h0c8c3: out <= 12'h000;
      20'h0c8c4: out <= 12'h000;
      20'h0c8c5: out <= 12'h000;
      20'h0c8c6: out <= 12'h000;
      20'h0c8c7: out <= 12'h000;
      20'h0c8c8: out <= 12'h000;
      20'h0c8c9: out <= 12'h000;
      20'h0c8ca: out <= 12'h000;
      20'h0c8cb: out <= 12'h000;
      20'h0c8cc: out <= 12'h000;
      20'h0c8cd: out <= 12'h000;
      20'h0c8ce: out <= 12'h000;
      20'h0c8cf: out <= 12'h000;
      20'h0c8d0: out <= 12'h000;
      20'h0c8d1: out <= 12'h000;
      20'h0c8d2: out <= 12'h000;
      20'h0c8d3: out <= 12'h000;
      20'h0c8d4: out <= 12'h000;
      20'h0c8d5: out <= 12'h000;
      20'h0c8d6: out <= 12'h000;
      20'h0c8d7: out <= 12'h000;
      20'h0c8d8: out <= 12'h000;
      20'h0c8d9: out <= 12'h000;
      20'h0c8da: out <= 12'h000;
      20'h0c8db: out <= 12'h000;
      20'h0c8dc: out <= 12'h000;
      20'h0c8dd: out <= 12'h000;
      20'h0c8de: out <= 12'h000;
      20'h0c8df: out <= 12'h000;
      20'h0c8e0: out <= 12'h000;
      20'h0c8e1: out <= 12'h000;
      20'h0c8e2: out <= 12'h000;
      20'h0c8e3: out <= 12'h000;
      20'h0c8e4: out <= 12'h000;
      20'h0c8e5: out <= 12'h000;
      20'h0c8e6: out <= 12'h000;
      20'h0c8e7: out <= 12'h000;
      20'h0c8e8: out <= 12'h000;
      20'h0c8e9: out <= 12'h000;
      20'h0c8ea: out <= 12'h000;
      20'h0c8eb: out <= 12'h000;
      20'h0c8ec: out <= 12'h000;
      20'h0c8ed: out <= 12'h000;
      20'h0c8ee: out <= 12'h000;
      20'h0c8ef: out <= 12'h000;
      20'h0c8f0: out <= 12'h000;
      20'h0c8f1: out <= 12'h000;
      20'h0c8f2: out <= 12'h000;
      20'h0c8f3: out <= 12'h000;
      20'h0c8f4: out <= 12'h000;
      20'h0c8f5: out <= 12'h000;
      20'h0c8f6: out <= 12'h000;
      20'h0c8f7: out <= 12'h000;
      20'h0c8f8: out <= 12'h000;
      20'h0c8f9: out <= 12'h000;
      20'h0c8fa: out <= 12'h000;
      20'h0c8fb: out <= 12'h000;
      20'h0c8fc: out <= 12'h603;
      20'h0c8fd: out <= 12'h603;
      20'h0c8fe: out <= 12'h603;
      20'h0c8ff: out <= 12'h603;
      20'h0c900: out <= 12'hb27;
      20'h0c901: out <= 12'hb27;
      20'h0c902: out <= 12'hb27;
      20'h0c903: out <= 12'hb27;
      20'h0c904: out <= 12'hb27;
      20'h0c905: out <= 12'hb27;
      20'h0c906: out <= 12'hb27;
      20'h0c907: out <= 12'hb27;
      20'h0c908: out <= 12'hb27;
      20'h0c909: out <= 12'hb27;
      20'h0c90a: out <= 12'hb27;
      20'h0c90b: out <= 12'hb27;
      20'h0c90c: out <= 12'hb27;
      20'h0c90d: out <= 12'hb27;
      20'h0c90e: out <= 12'hb27;
      20'h0c90f: out <= 12'hb27;
      20'h0c910: out <= 12'hb27;
      20'h0c911: out <= 12'hb27;
      20'h0c912: out <= 12'hb27;
      20'h0c913: out <= 12'hb27;
      20'h0c914: out <= 12'hb27;
      20'h0c915: out <= 12'hb27;
      20'h0c916: out <= 12'hb27;
      20'h0c917: out <= 12'hb27;
      20'h0c918: out <= 12'hb27;
      20'h0c919: out <= 12'hb27;
      20'h0c91a: out <= 12'hb27;
      20'h0c91b: out <= 12'hb27;
      20'h0c91c: out <= 12'hb27;
      20'h0c91d: out <= 12'hb27;
      20'h0c91e: out <= 12'hb27;
      20'h0c91f: out <= 12'hb27;
      20'h0c920: out <= 12'hb27;
      20'h0c921: out <= 12'hb27;
      20'h0c922: out <= 12'hb27;
      20'h0c923: out <= 12'hb27;
      20'h0c924: out <= 12'hb27;
      20'h0c925: out <= 12'hb27;
      20'h0c926: out <= 12'hb27;
      20'h0c927: out <= 12'hb27;
      20'h0c928: out <= 12'hb27;
      20'h0c929: out <= 12'hb27;
      20'h0c92a: out <= 12'hb27;
      20'h0c92b: out <= 12'hb27;
      20'h0c92c: out <= 12'hb27;
      20'h0c92d: out <= 12'hb27;
      20'h0c92e: out <= 12'hb27;
      20'h0c92f: out <= 12'hb27;
      20'h0c930: out <= 12'hb27;
      20'h0c931: out <= 12'hb27;
      20'h0c932: out <= 12'hb27;
      20'h0c933: out <= 12'hb27;
      20'h0c934: out <= 12'hb27;
      20'h0c935: out <= 12'hb27;
      20'h0c936: out <= 12'hb27;
      20'h0c937: out <= 12'hb27;
      20'h0c938: out <= 12'hb27;
      20'h0c939: out <= 12'hb27;
      20'h0c93a: out <= 12'hb27;
      20'h0c93b: out <= 12'hb27;
      20'h0c93c: out <= 12'hb27;
      20'h0c93d: out <= 12'hb27;
      20'h0c93e: out <= 12'hb27;
      20'h0c93f: out <= 12'hb27;
      20'h0c940: out <= 12'h088;
      20'h0c941: out <= 12'h088;
      20'h0c942: out <= 12'h088;
      20'h0c943: out <= 12'h088;
      20'h0c944: out <= 12'h088;
      20'h0c945: out <= 12'h088;
      20'h0c946: out <= 12'h088;
      20'h0c947: out <= 12'h088;
      20'h0c948: out <= 12'h088;
      20'h0c949: out <= 12'h088;
      20'h0c94a: out <= 12'h088;
      20'h0c94b: out <= 12'h088;
      20'h0c94c: out <= 12'h088;
      20'h0c94d: out <= 12'h088;
      20'h0c94e: out <= 12'h088;
      20'h0c94f: out <= 12'h088;
      20'h0c950: out <= 12'h088;
      20'h0c951: out <= 12'h088;
      20'h0c952: out <= 12'h088;
      20'h0c953: out <= 12'h088;
      20'h0c954: out <= 12'h088;
      20'h0c955: out <= 12'h088;
      20'h0c956: out <= 12'h088;
      20'h0c957: out <= 12'h088;
      20'h0c958: out <= 12'h088;
      20'h0c959: out <= 12'h088;
      20'h0c95a: out <= 12'h088;
      20'h0c95b: out <= 12'h088;
      20'h0c95c: out <= 12'h088;
      20'h0c95d: out <= 12'h088;
      20'h0c95e: out <= 12'h088;
      20'h0c95f: out <= 12'h088;
      20'h0c960: out <= 12'h088;
      20'h0c961: out <= 12'h088;
      20'h0c962: out <= 12'h088;
      20'h0c963: out <= 12'h088;
      20'h0c964: out <= 12'h088;
      20'h0c965: out <= 12'h088;
      20'h0c966: out <= 12'h088;
      20'h0c967: out <= 12'h088;
      20'h0c968: out <= 12'h088;
      20'h0c969: out <= 12'h088;
      20'h0c96a: out <= 12'h088;
      20'h0c96b: out <= 12'h088;
      20'h0c96c: out <= 12'h088;
      20'h0c96d: out <= 12'h088;
      20'h0c96e: out <= 12'h088;
      20'h0c96f: out <= 12'h088;
      20'h0c970: out <= 12'h088;
      20'h0c971: out <= 12'h088;
      20'h0c972: out <= 12'h088;
      20'h0c973: out <= 12'h088;
      20'h0c974: out <= 12'h088;
      20'h0c975: out <= 12'h088;
      20'h0c976: out <= 12'h088;
      20'h0c977: out <= 12'h088;
      20'h0c978: out <= 12'h088;
      20'h0c979: out <= 12'h088;
      20'h0c97a: out <= 12'h088;
      20'h0c97b: out <= 12'h088;
      20'h0c97c: out <= 12'h088;
      20'h0c97d: out <= 12'h088;
      20'h0c97e: out <= 12'h088;
      20'h0c97f: out <= 12'h088;
      20'h0c980: out <= 12'h088;
      20'h0c981: out <= 12'h088;
      20'h0c982: out <= 12'h088;
      20'h0c983: out <= 12'h088;
      20'h0c984: out <= 12'h088;
      20'h0c985: out <= 12'h088;
      20'h0c986: out <= 12'h088;
      20'h0c987: out <= 12'h088;
      20'h0c988: out <= 12'h088;
      20'h0c989: out <= 12'h088;
      20'h0c98a: out <= 12'h088;
      20'h0c98b: out <= 12'h088;
      20'h0c98c: out <= 12'h088;
      20'h0c98d: out <= 12'h088;
      20'h0c98e: out <= 12'h088;
      20'h0c98f: out <= 12'h088;
      20'h0c990: out <= 12'h088;
      20'h0c991: out <= 12'h088;
      20'h0c992: out <= 12'h088;
      20'h0c993: out <= 12'h088;
      20'h0c994: out <= 12'h088;
      20'h0c995: out <= 12'h088;
      20'h0c996: out <= 12'h088;
      20'h0c997: out <= 12'h088;
      20'h0c998: out <= 12'h088;
      20'h0c999: out <= 12'h088;
      20'h0c99a: out <= 12'h088;
      20'h0c99b: out <= 12'h088;
      20'h0c99c: out <= 12'h088;
      20'h0c99d: out <= 12'h088;
      20'h0c99e: out <= 12'h088;
      20'h0c99f: out <= 12'h088;
      20'h0c9a0: out <= 12'h088;
      20'h0c9a1: out <= 12'h088;
      20'h0c9a2: out <= 12'h088;
      20'h0c9a3: out <= 12'h088;
      20'h0c9a4: out <= 12'h088;
      20'h0c9a5: out <= 12'h088;
      20'h0c9a6: out <= 12'h088;
      20'h0c9a7: out <= 12'h088;
      20'h0c9a8: out <= 12'h088;
      20'h0c9a9: out <= 12'h222;
      20'h0c9aa: out <= 12'h222;
      20'h0c9ab: out <= 12'h222;
      20'h0c9ac: out <= 12'h222;
      20'h0c9ad: out <= 12'h222;
      20'h0c9ae: out <= 12'h222;
      20'h0c9af: out <= 12'h222;
      20'h0c9b0: out <= 12'h222;
      20'h0c9b1: out <= 12'h222;
      20'h0c9b2: out <= 12'h222;
      20'h0c9b3: out <= 12'h222;
      20'h0c9b4: out <= 12'h660;
      20'h0c9b5: out <= 12'h222;
      20'h0c9b6: out <= 12'h222;
      20'h0c9b7: out <= 12'h222;
      20'h0c9b8: out <= 12'h222;
      20'h0c9b9: out <= 12'h222;
      20'h0c9ba: out <= 12'h222;
      20'h0c9bb: out <= 12'h222;
      20'h0c9bc: out <= 12'h222;
      20'h0c9bd: out <= 12'h222;
      20'h0c9be: out <= 12'h222;
      20'h0c9bf: out <= 12'h222;
      20'h0c9c0: out <= 12'h603;
      20'h0c9c1: out <= 12'h603;
      20'h0c9c2: out <= 12'h603;
      20'h0c9c3: out <= 12'h603;
      20'h0c9c4: out <= 12'h603;
      20'h0c9c5: out <= 12'h603;
      20'h0c9c6: out <= 12'h603;
      20'h0c9c7: out <= 12'h603;
      20'h0c9c8: out <= 12'h603;
      20'h0c9c9: out <= 12'h603;
      20'h0c9ca: out <= 12'h603;
      20'h0c9cb: out <= 12'h603;
      20'h0c9cc: out <= 12'h603;
      20'h0c9cd: out <= 12'h603;
      20'h0c9ce: out <= 12'h603;
      20'h0c9cf: out <= 12'h603;
      20'h0c9d0: out <= 12'h603;
      20'h0c9d1: out <= 12'h603;
      20'h0c9d2: out <= 12'h603;
      20'h0c9d3: out <= 12'h603;
      20'h0c9d4: out <= 12'h603;
      20'h0c9d5: out <= 12'h603;
      20'h0c9d6: out <= 12'h603;
      20'h0c9d7: out <= 12'h603;
      20'h0c9d8: out <= 12'h603;
      20'h0c9d9: out <= 12'h603;
      20'h0c9da: out <= 12'h603;
      20'h0c9db: out <= 12'h603;
      20'h0c9dc: out <= 12'h603;
      20'h0c9dd: out <= 12'h603;
      20'h0c9de: out <= 12'h603;
      20'h0c9df: out <= 12'h603;
      20'h0c9e0: out <= 12'h603;
      20'h0c9e1: out <= 12'h603;
      20'h0c9e2: out <= 12'h603;
      20'h0c9e3: out <= 12'h603;
      20'h0c9e4: out <= 12'h603;
      20'h0c9e5: out <= 12'h603;
      20'h0c9e6: out <= 12'h603;
      20'h0c9e7: out <= 12'h603;
      20'h0c9e8: out <= 12'h603;
      20'h0c9e9: out <= 12'h603;
      20'h0c9ea: out <= 12'h603;
      20'h0c9eb: out <= 12'h603;
      20'h0c9ec: out <= 12'h603;
      20'h0c9ed: out <= 12'h603;
      20'h0c9ee: out <= 12'h603;
      20'h0c9ef: out <= 12'h603;
      20'h0c9f0: out <= 12'h603;
      20'h0c9f1: out <= 12'h603;
      20'h0c9f2: out <= 12'h603;
      20'h0c9f3: out <= 12'h603;
      20'h0c9f4: out <= 12'h603;
      20'h0c9f5: out <= 12'h603;
      20'h0c9f6: out <= 12'h603;
      20'h0c9f7: out <= 12'h603;
      20'h0c9f8: out <= 12'h603;
      20'h0c9f9: out <= 12'h603;
      20'h0c9fa: out <= 12'h603;
      20'h0c9fb: out <= 12'h603;
      20'h0c9fc: out <= 12'h603;
      20'h0c9fd: out <= 12'h603;
      20'h0c9fe: out <= 12'h603;
      20'h0c9ff: out <= 12'h603;
      20'h0ca00: out <= 12'h603;
      20'h0ca01: out <= 12'h603;
      20'h0ca02: out <= 12'h603;
      20'h0ca03: out <= 12'h603;
      20'h0ca04: out <= 12'h603;
      20'h0ca05: out <= 12'h603;
      20'h0ca06: out <= 12'h603;
      20'h0ca07: out <= 12'h603;
      20'h0ca08: out <= 12'h603;
      20'h0ca09: out <= 12'h603;
      20'h0ca0a: out <= 12'h603;
      20'h0ca0b: out <= 12'h603;
      20'h0ca0c: out <= 12'h603;
      20'h0ca0d: out <= 12'h603;
      20'h0ca0e: out <= 12'h603;
      20'h0ca0f: out <= 12'h603;
      20'h0ca10: out <= 12'h603;
      20'h0ca11: out <= 12'h603;
      20'h0ca12: out <= 12'h603;
      20'h0ca13: out <= 12'h603;
      20'h0ca14: out <= 12'h603;
      20'h0ca15: out <= 12'h603;
      20'h0ca16: out <= 12'h603;
      20'h0ca17: out <= 12'h603;
      20'h0ca18: out <= 12'hee9;
      20'h0ca19: out <= 12'hee9;
      20'h0ca1a: out <= 12'hee9;
      20'h0ca1b: out <= 12'hee9;
      20'h0ca1c: out <= 12'hee9;
      20'h0ca1d: out <= 12'hee9;
      20'h0ca1e: out <= 12'hee9;
      20'h0ca1f: out <= 12'hb27;
      20'h0ca20: out <= 12'h000;
      20'h0ca21: out <= 12'h000;
      20'h0ca22: out <= 12'h000;
      20'h0ca23: out <= 12'h000;
      20'h0ca24: out <= 12'h000;
      20'h0ca25: out <= 12'h000;
      20'h0ca26: out <= 12'h000;
      20'h0ca27: out <= 12'h000;
      20'h0ca28: out <= 12'h000;
      20'h0ca29: out <= 12'h000;
      20'h0ca2a: out <= 12'h000;
      20'h0ca2b: out <= 12'h000;
      20'h0ca2c: out <= 12'h000;
      20'h0ca2d: out <= 12'h000;
      20'h0ca2e: out <= 12'h000;
      20'h0ca2f: out <= 12'h000;
      20'h0ca30: out <= 12'h000;
      20'h0ca31: out <= 12'h000;
      20'h0ca32: out <= 12'h000;
      20'h0ca33: out <= 12'h000;
      20'h0ca34: out <= 12'h000;
      20'h0ca35: out <= 12'h000;
      20'h0ca36: out <= 12'h000;
      20'h0ca37: out <= 12'h000;
      20'h0ca38: out <= 12'h000;
      20'h0ca39: out <= 12'h000;
      20'h0ca3a: out <= 12'h000;
      20'h0ca3b: out <= 12'h000;
      20'h0ca3c: out <= 12'h000;
      20'h0ca3d: out <= 12'h000;
      20'h0ca3e: out <= 12'h000;
      20'h0ca3f: out <= 12'h000;
      20'h0ca40: out <= 12'h000;
      20'h0ca41: out <= 12'h000;
      20'h0ca42: out <= 12'h000;
      20'h0ca43: out <= 12'h000;
      20'h0ca44: out <= 12'h000;
      20'h0ca45: out <= 12'h000;
      20'h0ca46: out <= 12'h000;
      20'h0ca47: out <= 12'h000;
      20'h0ca48: out <= 12'h000;
      20'h0ca49: out <= 12'h000;
      20'h0ca4a: out <= 12'h000;
      20'h0ca4b: out <= 12'h000;
      20'h0ca4c: out <= 12'h000;
      20'h0ca4d: out <= 12'h000;
      20'h0ca4e: out <= 12'h000;
      20'h0ca4f: out <= 12'h000;
      20'h0ca50: out <= 12'h000;
      20'h0ca51: out <= 12'h000;
      20'h0ca52: out <= 12'h000;
      20'h0ca53: out <= 12'h000;
      20'h0ca54: out <= 12'h000;
      20'h0ca55: out <= 12'h000;
      20'h0ca56: out <= 12'h000;
      20'h0ca57: out <= 12'h000;
      20'h0ca58: out <= 12'h088;
      20'h0ca59: out <= 12'h088;
      20'h0ca5a: out <= 12'h088;
      20'h0ca5b: out <= 12'h088;
      20'h0ca5c: out <= 12'h088;
      20'h0ca5d: out <= 12'h088;
      20'h0ca5e: out <= 12'h088;
      20'h0ca5f: out <= 12'h088;
      20'h0ca60: out <= 12'h088;
      20'h0ca61: out <= 12'h088;
      20'h0ca62: out <= 12'h088;
      20'h0ca63: out <= 12'h088;
      20'h0ca64: out <= 12'h088;
      20'h0ca65: out <= 12'h088;
      20'h0ca66: out <= 12'h088;
      20'h0ca67: out <= 12'h088;
      20'h0ca68: out <= 12'h088;
      20'h0ca69: out <= 12'h088;
      20'h0ca6a: out <= 12'h088;
      20'h0ca6b: out <= 12'h088;
      20'h0ca6c: out <= 12'h088;
      20'h0ca6d: out <= 12'h088;
      20'h0ca6e: out <= 12'h088;
      20'h0ca6f: out <= 12'h088;
      20'h0ca70: out <= 12'h088;
      20'h0ca71: out <= 12'h088;
      20'h0ca72: out <= 12'h088;
      20'h0ca73: out <= 12'h088;
      20'h0ca74: out <= 12'h088;
      20'h0ca75: out <= 12'h088;
      20'h0ca76: out <= 12'h088;
      20'h0ca77: out <= 12'h088;
      20'h0ca78: out <= 12'h088;
      20'h0ca79: out <= 12'h088;
      20'h0ca7a: out <= 12'h088;
      20'h0ca7b: out <= 12'h088;
      20'h0ca7c: out <= 12'h088;
      20'h0ca7d: out <= 12'h088;
      20'h0ca7e: out <= 12'h088;
      20'h0ca7f: out <= 12'h088;
      20'h0ca80: out <= 12'h088;
      20'h0ca81: out <= 12'h088;
      20'h0ca82: out <= 12'h088;
      20'h0ca83: out <= 12'h088;
      20'h0ca84: out <= 12'h088;
      20'h0ca85: out <= 12'h088;
      20'h0ca86: out <= 12'h088;
      20'h0ca87: out <= 12'h088;
      20'h0ca88: out <= 12'h088;
      20'h0ca89: out <= 12'h088;
      20'h0ca8a: out <= 12'h088;
      20'h0ca8b: out <= 12'h088;
      20'h0ca8c: out <= 12'h088;
      20'h0ca8d: out <= 12'h088;
      20'h0ca8e: out <= 12'h088;
      20'h0ca8f: out <= 12'h088;
      20'h0ca90: out <= 12'h088;
      20'h0ca91: out <= 12'h088;
      20'h0ca92: out <= 12'h088;
      20'h0ca93: out <= 12'h088;
      20'h0ca94: out <= 12'h088;
      20'h0ca95: out <= 12'h088;
      20'h0ca96: out <= 12'h088;
      20'h0ca97: out <= 12'h088;
      20'h0ca98: out <= 12'h088;
      20'h0ca99: out <= 12'h088;
      20'h0ca9a: out <= 12'h088;
      20'h0ca9b: out <= 12'h088;
      20'h0ca9c: out <= 12'h088;
      20'h0ca9d: out <= 12'h088;
      20'h0ca9e: out <= 12'h088;
      20'h0ca9f: out <= 12'h088;
      20'h0caa0: out <= 12'h088;
      20'h0caa1: out <= 12'h088;
      20'h0caa2: out <= 12'h088;
      20'h0caa3: out <= 12'h088;
      20'h0caa4: out <= 12'h088;
      20'h0caa5: out <= 12'h088;
      20'h0caa6: out <= 12'h088;
      20'h0caa7: out <= 12'h088;
      20'h0caa8: out <= 12'h088;
      20'h0caa9: out <= 12'h088;
      20'h0caaa: out <= 12'h088;
      20'h0caab: out <= 12'h088;
      20'h0caac: out <= 12'h088;
      20'h0caad: out <= 12'h088;
      20'h0caae: out <= 12'h088;
      20'h0caaf: out <= 12'h088;
      20'h0cab0: out <= 12'h088;
      20'h0cab1: out <= 12'h088;
      20'h0cab2: out <= 12'h088;
      20'h0cab3: out <= 12'h088;
      20'h0cab4: out <= 12'h088;
      20'h0cab5: out <= 12'h088;
      20'h0cab6: out <= 12'h088;
      20'h0cab7: out <= 12'h088;
      20'h0cab8: out <= 12'h088;
      20'h0cab9: out <= 12'h088;
      20'h0caba: out <= 12'h088;
      20'h0cabb: out <= 12'h088;
      20'h0cabc: out <= 12'h088;
      20'h0cabd: out <= 12'h088;
      20'h0cabe: out <= 12'h088;
      20'h0cabf: out <= 12'h088;
      20'h0cac0: out <= 12'h088;
      20'h0cac1: out <= 12'h222;
      20'h0cac2: out <= 12'h222;
      20'h0cac3: out <= 12'h222;
      20'h0cac4: out <= 12'h222;
      20'h0cac5: out <= 12'h222;
      20'h0cac6: out <= 12'h222;
      20'h0cac7: out <= 12'h222;
      20'h0cac8: out <= 12'h222;
      20'h0cac9: out <= 12'h222;
      20'h0caca: out <= 12'h222;
      20'h0cacb: out <= 12'h222;
      20'h0cacc: out <= 12'h222;
      20'h0cacd: out <= 12'h222;
      20'h0cace: out <= 12'h222;
      20'h0cacf: out <= 12'h222;
      20'h0cad0: out <= 12'h222;
      20'h0cad1: out <= 12'h222;
      20'h0cad2: out <= 12'h222;
      20'h0cad3: out <= 12'h222;
      20'h0cad4: out <= 12'h222;
      20'h0cad5: out <= 12'h222;
      20'h0cad6: out <= 12'h222;
      20'h0cad7: out <= 12'h222;
      20'h0cad8: out <= 12'h603;
      20'h0cad9: out <= 12'h603;
      20'h0cada: out <= 12'h603;
      20'h0cadb: out <= 12'h603;
      20'h0cadc: out <= 12'h603;
      20'h0cadd: out <= 12'h603;
      20'h0cade: out <= 12'h603;
      20'h0cadf: out <= 12'h603;
      20'h0cae0: out <= 12'h603;
      20'h0cae1: out <= 12'h603;
      20'h0cae2: out <= 12'h603;
      20'h0cae3: out <= 12'h603;
      20'h0cae4: out <= 12'h603;
      20'h0cae5: out <= 12'h603;
      20'h0cae6: out <= 12'h603;
      20'h0cae7: out <= 12'h603;
      20'h0cae8: out <= 12'h603;
      20'h0cae9: out <= 12'h603;
      20'h0caea: out <= 12'h603;
      20'h0caeb: out <= 12'h603;
      20'h0caec: out <= 12'h603;
      20'h0caed: out <= 12'h603;
      20'h0caee: out <= 12'h603;
      20'h0caef: out <= 12'h603;
      20'h0caf0: out <= 12'h603;
      20'h0caf1: out <= 12'h603;
      20'h0caf2: out <= 12'h603;
      20'h0caf3: out <= 12'h603;
      20'h0caf4: out <= 12'h603;
      20'h0caf5: out <= 12'h603;
      20'h0caf6: out <= 12'h603;
      20'h0caf7: out <= 12'h603;
      20'h0caf8: out <= 12'h603;
      20'h0caf9: out <= 12'h603;
      20'h0cafa: out <= 12'h603;
      20'h0cafb: out <= 12'h603;
      20'h0cafc: out <= 12'h603;
      20'h0cafd: out <= 12'h603;
      20'h0cafe: out <= 12'h603;
      20'h0caff: out <= 12'h603;
      20'h0cb00: out <= 12'h603;
      20'h0cb01: out <= 12'h603;
      20'h0cb02: out <= 12'h603;
      20'h0cb03: out <= 12'h603;
      20'h0cb04: out <= 12'h603;
      20'h0cb05: out <= 12'h603;
      20'h0cb06: out <= 12'h603;
      20'h0cb07: out <= 12'h603;
      20'h0cb08: out <= 12'h603;
      20'h0cb09: out <= 12'h603;
      20'h0cb0a: out <= 12'h603;
      20'h0cb0b: out <= 12'h603;
      20'h0cb0c: out <= 12'h603;
      20'h0cb0d: out <= 12'h603;
      20'h0cb0e: out <= 12'h603;
      20'h0cb0f: out <= 12'h603;
      20'h0cb10: out <= 12'h603;
      20'h0cb11: out <= 12'h603;
      20'h0cb12: out <= 12'h603;
      20'h0cb13: out <= 12'h603;
      20'h0cb14: out <= 12'h603;
      20'h0cb15: out <= 12'h603;
      20'h0cb16: out <= 12'h603;
      20'h0cb17: out <= 12'h603;
      20'h0cb18: out <= 12'h603;
      20'h0cb19: out <= 12'h603;
      20'h0cb1a: out <= 12'h603;
      20'h0cb1b: out <= 12'h603;
      20'h0cb1c: out <= 12'h603;
      20'h0cb1d: out <= 12'h603;
      20'h0cb1e: out <= 12'h603;
      20'h0cb1f: out <= 12'h603;
      20'h0cb20: out <= 12'h603;
      20'h0cb21: out <= 12'h603;
      20'h0cb22: out <= 12'h603;
      20'h0cb23: out <= 12'h603;
      20'h0cb24: out <= 12'h603;
      20'h0cb25: out <= 12'h603;
      20'h0cb26: out <= 12'h603;
      20'h0cb27: out <= 12'h603;
      20'h0cb28: out <= 12'h603;
      20'h0cb29: out <= 12'h603;
      20'h0cb2a: out <= 12'h603;
      20'h0cb2b: out <= 12'h603;
      20'h0cb2c: out <= 12'h603;
      20'h0cb2d: out <= 12'h603;
      20'h0cb2e: out <= 12'h603;
      20'h0cb2f: out <= 12'h603;
      20'h0cb30: out <= 12'hee9;
      20'h0cb31: out <= 12'hf87;
      20'h0cb32: out <= 12'hf87;
      20'h0cb33: out <= 12'hf87;
      20'h0cb34: out <= 12'hf87;
      20'h0cb35: out <= 12'hf87;
      20'h0cb36: out <= 12'hf87;
      20'h0cb37: out <= 12'hb27;
      20'h0cb38: out <= 12'h000;
      20'h0cb39: out <= 12'h000;
      20'h0cb3a: out <= 12'h000;
      20'h0cb3b: out <= 12'h000;
      20'h0cb3c: out <= 12'h000;
      20'h0cb3d: out <= 12'h000;
      20'h0cb3e: out <= 12'h000;
      20'h0cb3f: out <= 12'h000;
      20'h0cb40: out <= 12'h000;
      20'h0cb41: out <= 12'h000;
      20'h0cb42: out <= 12'h000;
      20'h0cb43: out <= 12'h000;
      20'h0cb44: out <= 12'h000;
      20'h0cb45: out <= 12'h000;
      20'h0cb46: out <= 12'h000;
      20'h0cb47: out <= 12'h000;
      20'h0cb48: out <= 12'h000;
      20'h0cb49: out <= 12'h000;
      20'h0cb4a: out <= 12'h000;
      20'h0cb4b: out <= 12'h000;
      20'h0cb4c: out <= 12'h000;
      20'h0cb4d: out <= 12'h000;
      20'h0cb4e: out <= 12'h000;
      20'h0cb4f: out <= 12'h000;
      20'h0cb50: out <= 12'h000;
      20'h0cb51: out <= 12'h000;
      20'h0cb52: out <= 12'h000;
      20'h0cb53: out <= 12'h000;
      20'h0cb54: out <= 12'h000;
      20'h0cb55: out <= 12'h000;
      20'h0cb56: out <= 12'h000;
      20'h0cb57: out <= 12'h000;
      20'h0cb58: out <= 12'h000;
      20'h0cb59: out <= 12'h000;
      20'h0cb5a: out <= 12'h000;
      20'h0cb5b: out <= 12'h000;
      20'h0cb5c: out <= 12'h000;
      20'h0cb5d: out <= 12'h000;
      20'h0cb5e: out <= 12'h000;
      20'h0cb5f: out <= 12'h000;
      20'h0cb60: out <= 12'h000;
      20'h0cb61: out <= 12'h000;
      20'h0cb62: out <= 12'h000;
      20'h0cb63: out <= 12'h000;
      20'h0cb64: out <= 12'h000;
      20'h0cb65: out <= 12'h000;
      20'h0cb66: out <= 12'h000;
      20'h0cb67: out <= 12'h000;
      20'h0cb68: out <= 12'h000;
      20'h0cb69: out <= 12'h000;
      20'h0cb6a: out <= 12'h000;
      20'h0cb6b: out <= 12'h000;
      20'h0cb6c: out <= 12'h000;
      20'h0cb6d: out <= 12'h000;
      20'h0cb6e: out <= 12'h000;
      20'h0cb6f: out <= 12'h000;
      20'h0cb70: out <= 12'h088;
      20'h0cb71: out <= 12'h088;
      20'h0cb72: out <= 12'h088;
      20'h0cb73: out <= 12'h088;
      20'h0cb74: out <= 12'h088;
      20'h0cb75: out <= 12'h088;
      20'h0cb76: out <= 12'h088;
      20'h0cb77: out <= 12'h088;
      20'h0cb78: out <= 12'h088;
      20'h0cb79: out <= 12'h088;
      20'h0cb7a: out <= 12'h088;
      20'h0cb7b: out <= 12'h088;
      20'h0cb7c: out <= 12'h088;
      20'h0cb7d: out <= 12'h088;
      20'h0cb7e: out <= 12'h088;
      20'h0cb7f: out <= 12'h088;
      20'h0cb80: out <= 12'h088;
      20'h0cb81: out <= 12'h088;
      20'h0cb82: out <= 12'h088;
      20'h0cb83: out <= 12'h088;
      20'h0cb84: out <= 12'h088;
      20'h0cb85: out <= 12'h088;
      20'h0cb86: out <= 12'h088;
      20'h0cb87: out <= 12'h088;
      20'h0cb88: out <= 12'h088;
      20'h0cb89: out <= 12'h088;
      20'h0cb8a: out <= 12'h088;
      20'h0cb8b: out <= 12'h088;
      20'h0cb8c: out <= 12'h088;
      20'h0cb8d: out <= 12'h088;
      20'h0cb8e: out <= 12'h088;
      20'h0cb8f: out <= 12'h088;
      20'h0cb90: out <= 12'h088;
      20'h0cb91: out <= 12'h088;
      20'h0cb92: out <= 12'h088;
      20'h0cb93: out <= 12'h088;
      20'h0cb94: out <= 12'h088;
      20'h0cb95: out <= 12'h088;
      20'h0cb96: out <= 12'h088;
      20'h0cb97: out <= 12'h088;
      20'h0cb98: out <= 12'h088;
      20'h0cb99: out <= 12'h088;
      20'h0cb9a: out <= 12'h088;
      20'h0cb9b: out <= 12'h088;
      20'h0cb9c: out <= 12'h088;
      20'h0cb9d: out <= 12'h088;
      20'h0cb9e: out <= 12'h088;
      20'h0cb9f: out <= 12'h088;
      20'h0cba0: out <= 12'h088;
      20'h0cba1: out <= 12'h088;
      20'h0cba2: out <= 12'h088;
      20'h0cba3: out <= 12'h088;
      20'h0cba4: out <= 12'h088;
      20'h0cba5: out <= 12'h088;
      20'h0cba6: out <= 12'h088;
      20'h0cba7: out <= 12'h088;
      20'h0cba8: out <= 12'h088;
      20'h0cba9: out <= 12'h088;
      20'h0cbaa: out <= 12'h088;
      20'h0cbab: out <= 12'h088;
      20'h0cbac: out <= 12'h088;
      20'h0cbad: out <= 12'h088;
      20'h0cbae: out <= 12'h088;
      20'h0cbaf: out <= 12'h088;
      20'h0cbb0: out <= 12'h088;
      20'h0cbb1: out <= 12'h088;
      20'h0cbb2: out <= 12'h088;
      20'h0cbb3: out <= 12'h088;
      20'h0cbb4: out <= 12'h088;
      20'h0cbb5: out <= 12'h088;
      20'h0cbb6: out <= 12'h088;
      20'h0cbb7: out <= 12'h088;
      20'h0cbb8: out <= 12'h088;
      20'h0cbb9: out <= 12'h088;
      20'h0cbba: out <= 12'h088;
      20'h0cbbb: out <= 12'h088;
      20'h0cbbc: out <= 12'h088;
      20'h0cbbd: out <= 12'h088;
      20'h0cbbe: out <= 12'h088;
      20'h0cbbf: out <= 12'h088;
      20'h0cbc0: out <= 12'h088;
      20'h0cbc1: out <= 12'h088;
      20'h0cbc2: out <= 12'h088;
      20'h0cbc3: out <= 12'h088;
      20'h0cbc4: out <= 12'h088;
      20'h0cbc5: out <= 12'h088;
      20'h0cbc6: out <= 12'h088;
      20'h0cbc7: out <= 12'h088;
      20'h0cbc8: out <= 12'h088;
      20'h0cbc9: out <= 12'h088;
      20'h0cbca: out <= 12'h088;
      20'h0cbcb: out <= 12'h088;
      20'h0cbcc: out <= 12'h088;
      20'h0cbcd: out <= 12'h088;
      20'h0cbce: out <= 12'h088;
      20'h0cbcf: out <= 12'h088;
      20'h0cbd0: out <= 12'h088;
      20'h0cbd1: out <= 12'h088;
      20'h0cbd2: out <= 12'h088;
      20'h0cbd3: out <= 12'h088;
      20'h0cbd4: out <= 12'h088;
      20'h0cbd5: out <= 12'h088;
      20'h0cbd6: out <= 12'h088;
      20'h0cbd7: out <= 12'h088;
      20'h0cbd8: out <= 12'h088;
      20'h0cbd9: out <= 12'h222;
      20'h0cbda: out <= 12'h222;
      20'h0cbdb: out <= 12'h222;
      20'h0cbdc: out <= 12'h222;
      20'h0cbdd: out <= 12'h222;
      20'h0cbde: out <= 12'h222;
      20'h0cbdf: out <= 12'h222;
      20'h0cbe0: out <= 12'h222;
      20'h0cbe1: out <= 12'h222;
      20'h0cbe2: out <= 12'h222;
      20'h0cbe3: out <= 12'h222;
      20'h0cbe4: out <= 12'h222;
      20'h0cbe5: out <= 12'h222;
      20'h0cbe6: out <= 12'h222;
      20'h0cbe7: out <= 12'h222;
      20'h0cbe8: out <= 12'h222;
      20'h0cbe9: out <= 12'h222;
      20'h0cbea: out <= 12'h222;
      20'h0cbeb: out <= 12'h222;
      20'h0cbec: out <= 12'h222;
      20'h0cbed: out <= 12'h222;
      20'h0cbee: out <= 12'h222;
      20'h0cbef: out <= 12'h222;
      20'h0cbf0: out <= 12'h603;
      20'h0cbf1: out <= 12'h603;
      20'h0cbf2: out <= 12'h603;
      20'h0cbf3: out <= 12'h603;
      20'h0cbf4: out <= 12'h603;
      20'h0cbf5: out <= 12'h603;
      20'h0cbf6: out <= 12'h603;
      20'h0cbf7: out <= 12'h603;
      20'h0cbf8: out <= 12'h603;
      20'h0cbf9: out <= 12'h603;
      20'h0cbfa: out <= 12'h603;
      20'h0cbfb: out <= 12'h603;
      20'h0cbfc: out <= 12'h603;
      20'h0cbfd: out <= 12'h603;
      20'h0cbfe: out <= 12'h603;
      20'h0cbff: out <= 12'h603;
      20'h0cc00: out <= 12'h603;
      20'h0cc01: out <= 12'h603;
      20'h0cc02: out <= 12'h603;
      20'h0cc03: out <= 12'h603;
      20'h0cc04: out <= 12'h603;
      20'h0cc05: out <= 12'h603;
      20'h0cc06: out <= 12'h603;
      20'h0cc07: out <= 12'h603;
      20'h0cc08: out <= 12'h603;
      20'h0cc09: out <= 12'h603;
      20'h0cc0a: out <= 12'h603;
      20'h0cc0b: out <= 12'h603;
      20'h0cc0c: out <= 12'h603;
      20'h0cc0d: out <= 12'h603;
      20'h0cc0e: out <= 12'h603;
      20'h0cc0f: out <= 12'h603;
      20'h0cc10: out <= 12'h603;
      20'h0cc11: out <= 12'h603;
      20'h0cc12: out <= 12'h603;
      20'h0cc13: out <= 12'h603;
      20'h0cc14: out <= 12'h603;
      20'h0cc15: out <= 12'h603;
      20'h0cc16: out <= 12'h603;
      20'h0cc17: out <= 12'h603;
      20'h0cc18: out <= 12'h603;
      20'h0cc19: out <= 12'h603;
      20'h0cc1a: out <= 12'h603;
      20'h0cc1b: out <= 12'h603;
      20'h0cc1c: out <= 12'h603;
      20'h0cc1d: out <= 12'h603;
      20'h0cc1e: out <= 12'h603;
      20'h0cc1f: out <= 12'h603;
      20'h0cc20: out <= 12'h603;
      20'h0cc21: out <= 12'h603;
      20'h0cc22: out <= 12'h603;
      20'h0cc23: out <= 12'h603;
      20'h0cc24: out <= 12'h603;
      20'h0cc25: out <= 12'h603;
      20'h0cc26: out <= 12'h603;
      20'h0cc27: out <= 12'h603;
      20'h0cc28: out <= 12'h603;
      20'h0cc29: out <= 12'h603;
      20'h0cc2a: out <= 12'h603;
      20'h0cc2b: out <= 12'h603;
      20'h0cc2c: out <= 12'h603;
      20'h0cc2d: out <= 12'h603;
      20'h0cc2e: out <= 12'h603;
      20'h0cc2f: out <= 12'h603;
      20'h0cc30: out <= 12'h603;
      20'h0cc31: out <= 12'h603;
      20'h0cc32: out <= 12'h603;
      20'h0cc33: out <= 12'h603;
      20'h0cc34: out <= 12'h603;
      20'h0cc35: out <= 12'h603;
      20'h0cc36: out <= 12'h603;
      20'h0cc37: out <= 12'h603;
      20'h0cc38: out <= 12'h603;
      20'h0cc39: out <= 12'h603;
      20'h0cc3a: out <= 12'h603;
      20'h0cc3b: out <= 12'h603;
      20'h0cc3c: out <= 12'h603;
      20'h0cc3d: out <= 12'h603;
      20'h0cc3e: out <= 12'h603;
      20'h0cc3f: out <= 12'h603;
      20'h0cc40: out <= 12'h603;
      20'h0cc41: out <= 12'h603;
      20'h0cc42: out <= 12'h603;
      20'h0cc43: out <= 12'h603;
      20'h0cc44: out <= 12'h603;
      20'h0cc45: out <= 12'h603;
      20'h0cc46: out <= 12'h603;
      20'h0cc47: out <= 12'h603;
      20'h0cc48: out <= 12'hee9;
      20'h0cc49: out <= 12'hf87;
      20'h0cc4a: out <= 12'hee9;
      20'h0cc4b: out <= 12'hee9;
      20'h0cc4c: out <= 12'hee9;
      20'h0cc4d: out <= 12'hb27;
      20'h0cc4e: out <= 12'hf87;
      20'h0cc4f: out <= 12'hb27;
      20'h0cc50: out <= 12'h000;
      20'h0cc51: out <= 12'h000;
      20'h0cc52: out <= 12'h000;
      20'h0cc53: out <= 12'h000;
      20'h0cc54: out <= 12'h000;
      20'h0cc55: out <= 12'h000;
      20'h0cc56: out <= 12'h000;
      20'h0cc57: out <= 12'h000;
      20'h0cc58: out <= 12'h000;
      20'h0cc59: out <= 12'h000;
      20'h0cc5a: out <= 12'h000;
      20'h0cc5b: out <= 12'h000;
      20'h0cc5c: out <= 12'h000;
      20'h0cc5d: out <= 12'h000;
      20'h0cc5e: out <= 12'h000;
      20'h0cc5f: out <= 12'h000;
      20'h0cc60: out <= 12'h000;
      20'h0cc61: out <= 12'h000;
      20'h0cc62: out <= 12'h000;
      20'h0cc63: out <= 12'h000;
      20'h0cc64: out <= 12'h000;
      20'h0cc65: out <= 12'h000;
      20'h0cc66: out <= 12'h000;
      20'h0cc67: out <= 12'h000;
      20'h0cc68: out <= 12'h000;
      20'h0cc69: out <= 12'h000;
      20'h0cc6a: out <= 12'h000;
      20'h0cc6b: out <= 12'h000;
      20'h0cc6c: out <= 12'h000;
      20'h0cc6d: out <= 12'h000;
      20'h0cc6e: out <= 12'h000;
      20'h0cc6f: out <= 12'h000;
      20'h0cc70: out <= 12'h000;
      20'h0cc71: out <= 12'h000;
      20'h0cc72: out <= 12'h000;
      20'h0cc73: out <= 12'h000;
      20'h0cc74: out <= 12'h000;
      20'h0cc75: out <= 12'h000;
      20'h0cc76: out <= 12'h000;
      20'h0cc77: out <= 12'h000;
      20'h0cc78: out <= 12'h000;
      20'h0cc79: out <= 12'h000;
      20'h0cc7a: out <= 12'h000;
      20'h0cc7b: out <= 12'h000;
      20'h0cc7c: out <= 12'h000;
      20'h0cc7d: out <= 12'h000;
      20'h0cc7e: out <= 12'h000;
      20'h0cc7f: out <= 12'h000;
      20'h0cc80: out <= 12'h000;
      20'h0cc81: out <= 12'h000;
      20'h0cc82: out <= 12'h000;
      20'h0cc83: out <= 12'h000;
      20'h0cc84: out <= 12'h000;
      20'h0cc85: out <= 12'h000;
      20'h0cc86: out <= 12'h000;
      20'h0cc87: out <= 12'h000;
      20'h0cc88: out <= 12'h088;
      20'h0cc89: out <= 12'h088;
      20'h0cc8a: out <= 12'h088;
      20'h0cc8b: out <= 12'h088;
      20'h0cc8c: out <= 12'h088;
      20'h0cc8d: out <= 12'h088;
      20'h0cc8e: out <= 12'h088;
      20'h0cc8f: out <= 12'h088;
      20'h0cc90: out <= 12'h088;
      20'h0cc91: out <= 12'h088;
      20'h0cc92: out <= 12'h088;
      20'h0cc93: out <= 12'h088;
      20'h0cc94: out <= 12'h088;
      20'h0cc95: out <= 12'h088;
      20'h0cc96: out <= 12'h088;
      20'h0cc97: out <= 12'h088;
      20'h0cc98: out <= 12'h088;
      20'h0cc99: out <= 12'h088;
      20'h0cc9a: out <= 12'h088;
      20'h0cc9b: out <= 12'h088;
      20'h0cc9c: out <= 12'h088;
      20'h0cc9d: out <= 12'h088;
      20'h0cc9e: out <= 12'h088;
      20'h0cc9f: out <= 12'h088;
      20'h0cca0: out <= 12'h088;
      20'h0cca1: out <= 12'h088;
      20'h0cca2: out <= 12'h088;
      20'h0cca3: out <= 12'h088;
      20'h0cca4: out <= 12'h088;
      20'h0cca5: out <= 12'h088;
      20'h0cca6: out <= 12'h088;
      20'h0cca7: out <= 12'h088;
      20'h0cca8: out <= 12'h088;
      20'h0cca9: out <= 12'h088;
      20'h0ccaa: out <= 12'h088;
      20'h0ccab: out <= 12'h088;
      20'h0ccac: out <= 12'h088;
      20'h0ccad: out <= 12'h088;
      20'h0ccae: out <= 12'h088;
      20'h0ccaf: out <= 12'h088;
      20'h0ccb0: out <= 12'h088;
      20'h0ccb1: out <= 12'h088;
      20'h0ccb2: out <= 12'h088;
      20'h0ccb3: out <= 12'h088;
      20'h0ccb4: out <= 12'h088;
      20'h0ccb5: out <= 12'h088;
      20'h0ccb6: out <= 12'h088;
      20'h0ccb7: out <= 12'h088;
      20'h0ccb8: out <= 12'h088;
      20'h0ccb9: out <= 12'h088;
      20'h0ccba: out <= 12'h088;
      20'h0ccbb: out <= 12'h088;
      20'h0ccbc: out <= 12'h088;
      20'h0ccbd: out <= 12'h088;
      20'h0ccbe: out <= 12'h088;
      20'h0ccbf: out <= 12'h088;
      20'h0ccc0: out <= 12'h088;
      20'h0ccc1: out <= 12'h088;
      20'h0ccc2: out <= 12'h088;
      20'h0ccc3: out <= 12'h088;
      20'h0ccc4: out <= 12'h088;
      20'h0ccc5: out <= 12'h088;
      20'h0ccc6: out <= 12'h088;
      20'h0ccc7: out <= 12'h088;
      20'h0ccc8: out <= 12'h088;
      20'h0ccc9: out <= 12'h088;
      20'h0ccca: out <= 12'h088;
      20'h0cccb: out <= 12'h088;
      20'h0cccc: out <= 12'h088;
      20'h0cccd: out <= 12'h088;
      20'h0ccce: out <= 12'h088;
      20'h0cccf: out <= 12'h088;
      20'h0ccd0: out <= 12'h088;
      20'h0ccd1: out <= 12'h088;
      20'h0ccd2: out <= 12'h088;
      20'h0ccd3: out <= 12'h088;
      20'h0ccd4: out <= 12'h088;
      20'h0ccd5: out <= 12'h088;
      20'h0ccd6: out <= 12'h088;
      20'h0ccd7: out <= 12'h088;
      20'h0ccd8: out <= 12'h088;
      20'h0ccd9: out <= 12'h088;
      20'h0ccda: out <= 12'h088;
      20'h0ccdb: out <= 12'h088;
      20'h0ccdc: out <= 12'h088;
      20'h0ccdd: out <= 12'h088;
      20'h0ccde: out <= 12'h088;
      20'h0ccdf: out <= 12'h088;
      20'h0cce0: out <= 12'h088;
      20'h0cce1: out <= 12'h088;
      20'h0cce2: out <= 12'h088;
      20'h0cce3: out <= 12'h088;
      20'h0cce4: out <= 12'h088;
      20'h0cce5: out <= 12'h088;
      20'h0cce6: out <= 12'h088;
      20'h0cce7: out <= 12'h088;
      20'h0cce8: out <= 12'h088;
      20'h0cce9: out <= 12'h088;
      20'h0ccea: out <= 12'h088;
      20'h0cceb: out <= 12'h088;
      20'h0ccec: out <= 12'h088;
      20'h0cced: out <= 12'h088;
      20'h0ccee: out <= 12'h088;
      20'h0ccef: out <= 12'h088;
      20'h0ccf0: out <= 12'h088;
      20'h0ccf1: out <= 12'h222;
      20'h0ccf2: out <= 12'h222;
      20'h0ccf3: out <= 12'h222;
      20'h0ccf4: out <= 12'h222;
      20'h0ccf5: out <= 12'h222;
      20'h0ccf6: out <= 12'h222;
      20'h0ccf7: out <= 12'h222;
      20'h0ccf8: out <= 12'h222;
      20'h0ccf9: out <= 12'h222;
      20'h0ccfa: out <= 12'h222;
      20'h0ccfb: out <= 12'h222;
      20'h0ccfc: out <= 12'h222;
      20'h0ccfd: out <= 12'h222;
      20'h0ccfe: out <= 12'h222;
      20'h0ccff: out <= 12'h222;
      20'h0cd00: out <= 12'h222;
      20'h0cd01: out <= 12'h222;
      20'h0cd02: out <= 12'h222;
      20'h0cd03: out <= 12'h222;
      20'h0cd04: out <= 12'h222;
      20'h0cd05: out <= 12'h222;
      20'h0cd06: out <= 12'h222;
      20'h0cd07: out <= 12'h222;
      20'h0cd08: out <= 12'h603;
      20'h0cd09: out <= 12'h603;
      20'h0cd0a: out <= 12'h603;
      20'h0cd0b: out <= 12'h603;
      20'h0cd0c: out <= 12'h603;
      20'h0cd0d: out <= 12'h603;
      20'h0cd0e: out <= 12'h603;
      20'h0cd0f: out <= 12'h603;
      20'h0cd10: out <= 12'h603;
      20'h0cd11: out <= 12'h603;
      20'h0cd12: out <= 12'h603;
      20'h0cd13: out <= 12'h603;
      20'h0cd14: out <= 12'h603;
      20'h0cd15: out <= 12'h603;
      20'h0cd16: out <= 12'h603;
      20'h0cd17: out <= 12'h603;
      20'h0cd18: out <= 12'h603;
      20'h0cd19: out <= 12'h603;
      20'h0cd1a: out <= 12'h603;
      20'h0cd1b: out <= 12'h603;
      20'h0cd1c: out <= 12'h603;
      20'h0cd1d: out <= 12'h603;
      20'h0cd1e: out <= 12'h603;
      20'h0cd1f: out <= 12'h603;
      20'h0cd20: out <= 12'h603;
      20'h0cd21: out <= 12'h603;
      20'h0cd22: out <= 12'h603;
      20'h0cd23: out <= 12'h603;
      20'h0cd24: out <= 12'h603;
      20'h0cd25: out <= 12'h603;
      20'h0cd26: out <= 12'h603;
      20'h0cd27: out <= 12'h603;
      20'h0cd28: out <= 12'h603;
      20'h0cd29: out <= 12'h603;
      20'h0cd2a: out <= 12'h603;
      20'h0cd2b: out <= 12'h603;
      20'h0cd2c: out <= 12'h603;
      20'h0cd2d: out <= 12'h603;
      20'h0cd2e: out <= 12'h603;
      20'h0cd2f: out <= 12'h603;
      20'h0cd30: out <= 12'h603;
      20'h0cd31: out <= 12'h603;
      20'h0cd32: out <= 12'h603;
      20'h0cd33: out <= 12'h603;
      20'h0cd34: out <= 12'h603;
      20'h0cd35: out <= 12'h603;
      20'h0cd36: out <= 12'h603;
      20'h0cd37: out <= 12'h603;
      20'h0cd38: out <= 12'h603;
      20'h0cd39: out <= 12'h603;
      20'h0cd3a: out <= 12'h603;
      20'h0cd3b: out <= 12'h603;
      20'h0cd3c: out <= 12'h603;
      20'h0cd3d: out <= 12'h603;
      20'h0cd3e: out <= 12'h603;
      20'h0cd3f: out <= 12'h603;
      20'h0cd40: out <= 12'h603;
      20'h0cd41: out <= 12'h603;
      20'h0cd42: out <= 12'h603;
      20'h0cd43: out <= 12'h603;
      20'h0cd44: out <= 12'h603;
      20'h0cd45: out <= 12'h603;
      20'h0cd46: out <= 12'h603;
      20'h0cd47: out <= 12'h603;
      20'h0cd48: out <= 12'h603;
      20'h0cd49: out <= 12'h603;
      20'h0cd4a: out <= 12'h603;
      20'h0cd4b: out <= 12'h603;
      20'h0cd4c: out <= 12'h603;
      20'h0cd4d: out <= 12'h603;
      20'h0cd4e: out <= 12'h603;
      20'h0cd4f: out <= 12'h603;
      20'h0cd50: out <= 12'h603;
      20'h0cd51: out <= 12'h603;
      20'h0cd52: out <= 12'h603;
      20'h0cd53: out <= 12'h603;
      20'h0cd54: out <= 12'h603;
      20'h0cd55: out <= 12'h603;
      20'h0cd56: out <= 12'h603;
      20'h0cd57: out <= 12'h603;
      20'h0cd58: out <= 12'h603;
      20'h0cd59: out <= 12'h603;
      20'h0cd5a: out <= 12'h603;
      20'h0cd5b: out <= 12'h603;
      20'h0cd5c: out <= 12'h603;
      20'h0cd5d: out <= 12'h603;
      20'h0cd5e: out <= 12'h603;
      20'h0cd5f: out <= 12'h603;
      20'h0cd60: out <= 12'hee9;
      20'h0cd61: out <= 12'hf87;
      20'h0cd62: out <= 12'hee9;
      20'h0cd63: out <= 12'hf87;
      20'h0cd64: out <= 12'hf87;
      20'h0cd65: out <= 12'hb27;
      20'h0cd66: out <= 12'hf87;
      20'h0cd67: out <= 12'hb27;
      20'h0cd68: out <= 12'h000;
      20'h0cd69: out <= 12'h000;
      20'h0cd6a: out <= 12'h000;
      20'h0cd6b: out <= 12'h000;
      20'h0cd6c: out <= 12'h000;
      20'h0cd6d: out <= 12'h000;
      20'h0cd6e: out <= 12'h000;
      20'h0cd6f: out <= 12'h000;
      20'h0cd70: out <= 12'h000;
      20'h0cd71: out <= 12'h000;
      20'h0cd72: out <= 12'h000;
      20'h0cd73: out <= 12'h000;
      20'h0cd74: out <= 12'h000;
      20'h0cd75: out <= 12'h000;
      20'h0cd76: out <= 12'h000;
      20'h0cd77: out <= 12'h000;
      20'h0cd78: out <= 12'h000;
      20'h0cd79: out <= 12'h000;
      20'h0cd7a: out <= 12'h000;
      20'h0cd7b: out <= 12'h000;
      20'h0cd7c: out <= 12'h000;
      20'h0cd7d: out <= 12'h000;
      20'h0cd7e: out <= 12'h000;
      20'h0cd7f: out <= 12'h000;
      20'h0cd80: out <= 12'h000;
      20'h0cd81: out <= 12'h000;
      20'h0cd82: out <= 12'h000;
      20'h0cd83: out <= 12'h000;
      20'h0cd84: out <= 12'h000;
      20'h0cd85: out <= 12'h000;
      20'h0cd86: out <= 12'h000;
      20'h0cd87: out <= 12'h000;
      20'h0cd88: out <= 12'h000;
      20'h0cd89: out <= 12'h000;
      20'h0cd8a: out <= 12'h000;
      20'h0cd8b: out <= 12'h000;
      20'h0cd8c: out <= 12'h000;
      20'h0cd8d: out <= 12'h000;
      20'h0cd8e: out <= 12'h000;
      20'h0cd8f: out <= 12'h000;
      20'h0cd90: out <= 12'h000;
      20'h0cd91: out <= 12'h000;
      20'h0cd92: out <= 12'h000;
      20'h0cd93: out <= 12'h000;
      20'h0cd94: out <= 12'h000;
      20'h0cd95: out <= 12'h000;
      20'h0cd96: out <= 12'h000;
      20'h0cd97: out <= 12'h000;
      20'h0cd98: out <= 12'h000;
      20'h0cd99: out <= 12'h000;
      20'h0cd9a: out <= 12'h000;
      20'h0cd9b: out <= 12'h000;
      20'h0cd9c: out <= 12'h000;
      20'h0cd9d: out <= 12'h000;
      20'h0cd9e: out <= 12'h000;
      20'h0cd9f: out <= 12'h000;
      20'h0cda0: out <= 12'h088;
      20'h0cda1: out <= 12'h088;
      20'h0cda2: out <= 12'h088;
      20'h0cda3: out <= 12'h088;
      20'h0cda4: out <= 12'h088;
      20'h0cda5: out <= 12'h088;
      20'h0cda6: out <= 12'h088;
      20'h0cda7: out <= 12'h088;
      20'h0cda8: out <= 12'h088;
      20'h0cda9: out <= 12'h088;
      20'h0cdaa: out <= 12'h088;
      20'h0cdab: out <= 12'h088;
      20'h0cdac: out <= 12'h088;
      20'h0cdad: out <= 12'h088;
      20'h0cdae: out <= 12'h088;
      20'h0cdaf: out <= 12'h088;
      20'h0cdb0: out <= 12'h088;
      20'h0cdb1: out <= 12'h088;
      20'h0cdb2: out <= 12'h088;
      20'h0cdb3: out <= 12'h088;
      20'h0cdb4: out <= 12'h088;
      20'h0cdb5: out <= 12'h088;
      20'h0cdb6: out <= 12'h088;
      20'h0cdb7: out <= 12'h088;
      20'h0cdb8: out <= 12'h088;
      20'h0cdb9: out <= 12'h088;
      20'h0cdba: out <= 12'h088;
      20'h0cdbb: out <= 12'h088;
      20'h0cdbc: out <= 12'h088;
      20'h0cdbd: out <= 12'h088;
      20'h0cdbe: out <= 12'h088;
      20'h0cdbf: out <= 12'h088;
      20'h0cdc0: out <= 12'h088;
      20'h0cdc1: out <= 12'h088;
      20'h0cdc2: out <= 12'h088;
      20'h0cdc3: out <= 12'h088;
      20'h0cdc4: out <= 12'h088;
      20'h0cdc5: out <= 12'h088;
      20'h0cdc6: out <= 12'h088;
      20'h0cdc7: out <= 12'h088;
      20'h0cdc8: out <= 12'h088;
      20'h0cdc9: out <= 12'h088;
      20'h0cdca: out <= 12'h088;
      20'h0cdcb: out <= 12'h088;
      20'h0cdcc: out <= 12'h088;
      20'h0cdcd: out <= 12'h088;
      20'h0cdce: out <= 12'h088;
      20'h0cdcf: out <= 12'h088;
      20'h0cdd0: out <= 12'h088;
      20'h0cdd1: out <= 12'h088;
      20'h0cdd2: out <= 12'h088;
      20'h0cdd3: out <= 12'h088;
      20'h0cdd4: out <= 12'h088;
      20'h0cdd5: out <= 12'h088;
      20'h0cdd6: out <= 12'h088;
      20'h0cdd7: out <= 12'h088;
      20'h0cdd8: out <= 12'h088;
      20'h0cdd9: out <= 12'h088;
      20'h0cdda: out <= 12'h088;
      20'h0cddb: out <= 12'h088;
      20'h0cddc: out <= 12'h088;
      20'h0cddd: out <= 12'h088;
      20'h0cdde: out <= 12'h088;
      20'h0cddf: out <= 12'h088;
      20'h0cde0: out <= 12'h088;
      20'h0cde1: out <= 12'h088;
      20'h0cde2: out <= 12'h088;
      20'h0cde3: out <= 12'h088;
      20'h0cde4: out <= 12'h088;
      20'h0cde5: out <= 12'h088;
      20'h0cde6: out <= 12'h088;
      20'h0cde7: out <= 12'h088;
      20'h0cde8: out <= 12'h088;
      20'h0cde9: out <= 12'h088;
      20'h0cdea: out <= 12'h088;
      20'h0cdeb: out <= 12'h088;
      20'h0cdec: out <= 12'h088;
      20'h0cded: out <= 12'h088;
      20'h0cdee: out <= 12'h088;
      20'h0cdef: out <= 12'h088;
      20'h0cdf0: out <= 12'h088;
      20'h0cdf1: out <= 12'h088;
      20'h0cdf2: out <= 12'h088;
      20'h0cdf3: out <= 12'h088;
      20'h0cdf4: out <= 12'h088;
      20'h0cdf5: out <= 12'h088;
      20'h0cdf6: out <= 12'h088;
      20'h0cdf7: out <= 12'h088;
      20'h0cdf8: out <= 12'h088;
      20'h0cdf9: out <= 12'h088;
      20'h0cdfa: out <= 12'h088;
      20'h0cdfb: out <= 12'h088;
      20'h0cdfc: out <= 12'h088;
      20'h0cdfd: out <= 12'h088;
      20'h0cdfe: out <= 12'h088;
      20'h0cdff: out <= 12'h088;
      20'h0ce00: out <= 12'h088;
      20'h0ce01: out <= 12'h088;
      20'h0ce02: out <= 12'h088;
      20'h0ce03: out <= 12'h088;
      20'h0ce04: out <= 12'h088;
      20'h0ce05: out <= 12'h088;
      20'h0ce06: out <= 12'h088;
      20'h0ce07: out <= 12'h088;
      20'h0ce08: out <= 12'h088;
      20'h0ce09: out <= 12'h603;
      20'h0ce0a: out <= 12'h603;
      20'h0ce0b: out <= 12'h603;
      20'h0ce0c: out <= 12'h603;
      20'h0ce0d: out <= 12'h603;
      20'h0ce0e: out <= 12'h603;
      20'h0ce0f: out <= 12'h603;
      20'h0ce10: out <= 12'h603;
      20'h0ce11: out <= 12'h603;
      20'h0ce12: out <= 12'h603;
      20'h0ce13: out <= 12'h603;
      20'h0ce14: out <= 12'h603;
      20'h0ce15: out <= 12'h603;
      20'h0ce16: out <= 12'h603;
      20'h0ce17: out <= 12'h603;
      20'h0ce18: out <= 12'h603;
      20'h0ce19: out <= 12'h603;
      20'h0ce1a: out <= 12'h603;
      20'h0ce1b: out <= 12'h603;
      20'h0ce1c: out <= 12'h603;
      20'h0ce1d: out <= 12'h603;
      20'h0ce1e: out <= 12'h603;
      20'h0ce1f: out <= 12'h603;
      20'h0ce20: out <= 12'h603;
      20'h0ce21: out <= 12'h603;
      20'h0ce22: out <= 12'h603;
      20'h0ce23: out <= 12'h603;
      20'h0ce24: out <= 12'h603;
      20'h0ce25: out <= 12'h603;
      20'h0ce26: out <= 12'h603;
      20'h0ce27: out <= 12'h603;
      20'h0ce28: out <= 12'h603;
      20'h0ce29: out <= 12'h603;
      20'h0ce2a: out <= 12'h603;
      20'h0ce2b: out <= 12'h603;
      20'h0ce2c: out <= 12'h603;
      20'h0ce2d: out <= 12'h603;
      20'h0ce2e: out <= 12'h603;
      20'h0ce2f: out <= 12'h603;
      20'h0ce30: out <= 12'h603;
      20'h0ce31: out <= 12'h603;
      20'h0ce32: out <= 12'h603;
      20'h0ce33: out <= 12'h603;
      20'h0ce34: out <= 12'h603;
      20'h0ce35: out <= 12'h603;
      20'h0ce36: out <= 12'h603;
      20'h0ce37: out <= 12'h603;
      20'h0ce38: out <= 12'h603;
      20'h0ce39: out <= 12'h603;
      20'h0ce3a: out <= 12'h603;
      20'h0ce3b: out <= 12'h603;
      20'h0ce3c: out <= 12'h603;
      20'h0ce3d: out <= 12'h603;
      20'h0ce3e: out <= 12'h603;
      20'h0ce3f: out <= 12'h603;
      20'h0ce40: out <= 12'h603;
      20'h0ce41: out <= 12'h603;
      20'h0ce42: out <= 12'h603;
      20'h0ce43: out <= 12'h603;
      20'h0ce44: out <= 12'h603;
      20'h0ce45: out <= 12'h603;
      20'h0ce46: out <= 12'h603;
      20'h0ce47: out <= 12'h603;
      20'h0ce48: out <= 12'h603;
      20'h0ce49: out <= 12'h603;
      20'h0ce4a: out <= 12'h603;
      20'h0ce4b: out <= 12'h603;
      20'h0ce4c: out <= 12'h603;
      20'h0ce4d: out <= 12'h603;
      20'h0ce4e: out <= 12'h603;
      20'h0ce4f: out <= 12'h603;
      20'h0ce50: out <= 12'h603;
      20'h0ce51: out <= 12'h603;
      20'h0ce52: out <= 12'h603;
      20'h0ce53: out <= 12'h603;
      20'h0ce54: out <= 12'h603;
      20'h0ce55: out <= 12'h603;
      20'h0ce56: out <= 12'h603;
      20'h0ce57: out <= 12'h603;
      20'h0ce58: out <= 12'h603;
      20'h0ce59: out <= 12'h603;
      20'h0ce5a: out <= 12'h603;
      20'h0ce5b: out <= 12'h603;
      20'h0ce5c: out <= 12'h603;
      20'h0ce5d: out <= 12'h603;
      20'h0ce5e: out <= 12'h603;
      20'h0ce5f: out <= 12'h603;
      20'h0ce60: out <= 12'h603;
      20'h0ce61: out <= 12'h603;
      20'h0ce62: out <= 12'h603;
      20'h0ce63: out <= 12'h603;
      20'h0ce64: out <= 12'h603;
      20'h0ce65: out <= 12'h603;
      20'h0ce66: out <= 12'h603;
      20'h0ce67: out <= 12'h603;
      20'h0ce68: out <= 12'h603;
      20'h0ce69: out <= 12'h603;
      20'h0ce6a: out <= 12'h603;
      20'h0ce6b: out <= 12'h603;
      20'h0ce6c: out <= 12'h603;
      20'h0ce6d: out <= 12'h603;
      20'h0ce6e: out <= 12'h603;
      20'h0ce6f: out <= 12'h603;
      20'h0ce70: out <= 12'h603;
      20'h0ce71: out <= 12'h603;
      20'h0ce72: out <= 12'h603;
      20'h0ce73: out <= 12'h603;
      20'h0ce74: out <= 12'h603;
      20'h0ce75: out <= 12'h603;
      20'h0ce76: out <= 12'h603;
      20'h0ce77: out <= 12'h603;
      20'h0ce78: out <= 12'hee9;
      20'h0ce79: out <= 12'hf87;
      20'h0ce7a: out <= 12'hee9;
      20'h0ce7b: out <= 12'hf87;
      20'h0ce7c: out <= 12'hf87;
      20'h0ce7d: out <= 12'hb27;
      20'h0ce7e: out <= 12'hf87;
      20'h0ce7f: out <= 12'hb27;
      20'h0ce80: out <= 12'h000;
      20'h0ce81: out <= 12'h000;
      20'h0ce82: out <= 12'h000;
      20'h0ce83: out <= 12'h000;
      20'h0ce84: out <= 12'h000;
      20'h0ce85: out <= 12'h000;
      20'h0ce86: out <= 12'h000;
      20'h0ce87: out <= 12'h000;
      20'h0ce88: out <= 12'h000;
      20'h0ce89: out <= 12'h000;
      20'h0ce8a: out <= 12'h000;
      20'h0ce8b: out <= 12'h000;
      20'h0ce8c: out <= 12'h000;
      20'h0ce8d: out <= 12'h000;
      20'h0ce8e: out <= 12'h000;
      20'h0ce8f: out <= 12'h000;
      20'h0ce90: out <= 12'h000;
      20'h0ce91: out <= 12'h000;
      20'h0ce92: out <= 12'h000;
      20'h0ce93: out <= 12'h000;
      20'h0ce94: out <= 12'h000;
      20'h0ce95: out <= 12'h000;
      20'h0ce96: out <= 12'h000;
      20'h0ce97: out <= 12'h000;
      20'h0ce98: out <= 12'h000;
      20'h0ce99: out <= 12'h000;
      20'h0ce9a: out <= 12'h000;
      20'h0ce9b: out <= 12'h000;
      20'h0ce9c: out <= 12'h000;
      20'h0ce9d: out <= 12'h000;
      20'h0ce9e: out <= 12'h000;
      20'h0ce9f: out <= 12'h000;
      20'h0cea0: out <= 12'h000;
      20'h0cea1: out <= 12'h000;
      20'h0cea2: out <= 12'h000;
      20'h0cea3: out <= 12'h000;
      20'h0cea4: out <= 12'h000;
      20'h0cea5: out <= 12'h000;
      20'h0cea6: out <= 12'h000;
      20'h0cea7: out <= 12'h000;
      20'h0cea8: out <= 12'h000;
      20'h0cea9: out <= 12'h000;
      20'h0ceaa: out <= 12'h000;
      20'h0ceab: out <= 12'h000;
      20'h0ceac: out <= 12'h000;
      20'h0cead: out <= 12'h000;
      20'h0ceae: out <= 12'h000;
      20'h0ceaf: out <= 12'h000;
      20'h0ceb0: out <= 12'h000;
      20'h0ceb1: out <= 12'h000;
      20'h0ceb2: out <= 12'h000;
      20'h0ceb3: out <= 12'h000;
      20'h0ceb4: out <= 12'h000;
      20'h0ceb5: out <= 12'h000;
      20'h0ceb6: out <= 12'h000;
      20'h0ceb7: out <= 12'h000;
      20'h0ceb8: out <= 12'h088;
      20'h0ceb9: out <= 12'h088;
      20'h0ceba: out <= 12'h088;
      20'h0cebb: out <= 12'h088;
      20'h0cebc: out <= 12'h088;
      20'h0cebd: out <= 12'h088;
      20'h0cebe: out <= 12'h088;
      20'h0cebf: out <= 12'h088;
      20'h0cec0: out <= 12'h088;
      20'h0cec1: out <= 12'h088;
      20'h0cec2: out <= 12'h088;
      20'h0cec3: out <= 12'h088;
      20'h0cec4: out <= 12'h088;
      20'h0cec5: out <= 12'h088;
      20'h0cec6: out <= 12'h088;
      20'h0cec7: out <= 12'h088;
      20'h0cec8: out <= 12'h088;
      20'h0cec9: out <= 12'h088;
      20'h0ceca: out <= 12'h088;
      20'h0cecb: out <= 12'h088;
      20'h0cecc: out <= 12'h088;
      20'h0cecd: out <= 12'h088;
      20'h0cece: out <= 12'h088;
      20'h0cecf: out <= 12'h088;
      20'h0ced0: out <= 12'h088;
      20'h0ced1: out <= 12'h088;
      20'h0ced2: out <= 12'h088;
      20'h0ced3: out <= 12'h088;
      20'h0ced4: out <= 12'h088;
      20'h0ced5: out <= 12'h088;
      20'h0ced6: out <= 12'h088;
      20'h0ced7: out <= 12'h088;
      20'h0ced8: out <= 12'h088;
      20'h0ced9: out <= 12'h088;
      20'h0ceda: out <= 12'h088;
      20'h0cedb: out <= 12'h088;
      20'h0cedc: out <= 12'h088;
      20'h0cedd: out <= 12'h088;
      20'h0cede: out <= 12'h088;
      20'h0cedf: out <= 12'h088;
      20'h0cee0: out <= 12'h088;
      20'h0cee1: out <= 12'h088;
      20'h0cee2: out <= 12'h088;
      20'h0cee3: out <= 12'h088;
      20'h0cee4: out <= 12'h088;
      20'h0cee5: out <= 12'h088;
      20'h0cee6: out <= 12'h088;
      20'h0cee7: out <= 12'h088;
      20'h0cee8: out <= 12'h088;
      20'h0cee9: out <= 12'h088;
      20'h0ceea: out <= 12'h088;
      20'h0ceeb: out <= 12'h088;
      20'h0ceec: out <= 12'h088;
      20'h0ceed: out <= 12'h088;
      20'h0ceee: out <= 12'h088;
      20'h0ceef: out <= 12'h088;
      20'h0cef0: out <= 12'h088;
      20'h0cef1: out <= 12'h088;
      20'h0cef2: out <= 12'h088;
      20'h0cef3: out <= 12'h088;
      20'h0cef4: out <= 12'h088;
      20'h0cef5: out <= 12'h088;
      20'h0cef6: out <= 12'h088;
      20'h0cef7: out <= 12'h088;
      20'h0cef8: out <= 12'h088;
      20'h0cef9: out <= 12'h088;
      20'h0cefa: out <= 12'h088;
      20'h0cefb: out <= 12'h088;
      20'h0cefc: out <= 12'h088;
      20'h0cefd: out <= 12'h088;
      20'h0cefe: out <= 12'h088;
      20'h0ceff: out <= 12'h088;
      20'h0cf00: out <= 12'h088;
      20'h0cf01: out <= 12'h088;
      20'h0cf02: out <= 12'h088;
      20'h0cf03: out <= 12'h088;
      20'h0cf04: out <= 12'h088;
      20'h0cf05: out <= 12'h088;
      20'h0cf06: out <= 12'h088;
      20'h0cf07: out <= 12'h088;
      20'h0cf08: out <= 12'h088;
      20'h0cf09: out <= 12'h088;
      20'h0cf0a: out <= 12'h088;
      20'h0cf0b: out <= 12'h088;
      20'h0cf0c: out <= 12'h088;
      20'h0cf0d: out <= 12'h088;
      20'h0cf0e: out <= 12'h088;
      20'h0cf0f: out <= 12'h088;
      20'h0cf10: out <= 12'h088;
      20'h0cf11: out <= 12'h088;
      20'h0cf12: out <= 12'h088;
      20'h0cf13: out <= 12'h088;
      20'h0cf14: out <= 12'h088;
      20'h0cf15: out <= 12'h088;
      20'h0cf16: out <= 12'h088;
      20'h0cf17: out <= 12'h088;
      20'h0cf18: out <= 12'h088;
      20'h0cf19: out <= 12'h088;
      20'h0cf1a: out <= 12'h088;
      20'h0cf1b: out <= 12'h088;
      20'h0cf1c: out <= 12'h088;
      20'h0cf1d: out <= 12'h088;
      20'h0cf1e: out <= 12'h088;
      20'h0cf1f: out <= 12'h088;
      20'h0cf20: out <= 12'h088;
      20'h0cf21: out <= 12'h603;
      20'h0cf22: out <= 12'h603;
      20'h0cf23: out <= 12'h603;
      20'h0cf24: out <= 12'h603;
      20'h0cf25: out <= 12'h603;
      20'h0cf26: out <= 12'h603;
      20'h0cf27: out <= 12'h603;
      20'h0cf28: out <= 12'h603;
      20'h0cf29: out <= 12'h603;
      20'h0cf2a: out <= 12'h603;
      20'h0cf2b: out <= 12'h603;
      20'h0cf2c: out <= 12'h603;
      20'h0cf2d: out <= 12'h603;
      20'h0cf2e: out <= 12'h603;
      20'h0cf2f: out <= 12'h603;
      20'h0cf30: out <= 12'h603;
      20'h0cf31: out <= 12'h603;
      20'h0cf32: out <= 12'h603;
      20'h0cf33: out <= 12'h603;
      20'h0cf34: out <= 12'h603;
      20'h0cf35: out <= 12'h603;
      20'h0cf36: out <= 12'h603;
      20'h0cf37: out <= 12'h603;
      20'h0cf38: out <= 12'h603;
      20'h0cf39: out <= 12'h603;
      20'h0cf3a: out <= 12'h603;
      20'h0cf3b: out <= 12'h603;
      20'h0cf3c: out <= 12'h603;
      20'h0cf3d: out <= 12'h603;
      20'h0cf3e: out <= 12'h603;
      20'h0cf3f: out <= 12'h603;
      20'h0cf40: out <= 12'h603;
      20'h0cf41: out <= 12'h603;
      20'h0cf42: out <= 12'h603;
      20'h0cf43: out <= 12'h603;
      20'h0cf44: out <= 12'h603;
      20'h0cf45: out <= 12'h603;
      20'h0cf46: out <= 12'h603;
      20'h0cf47: out <= 12'h603;
      20'h0cf48: out <= 12'h603;
      20'h0cf49: out <= 12'h603;
      20'h0cf4a: out <= 12'h603;
      20'h0cf4b: out <= 12'h603;
      20'h0cf4c: out <= 12'h603;
      20'h0cf4d: out <= 12'h603;
      20'h0cf4e: out <= 12'h603;
      20'h0cf4f: out <= 12'h603;
      20'h0cf50: out <= 12'h603;
      20'h0cf51: out <= 12'h603;
      20'h0cf52: out <= 12'h603;
      20'h0cf53: out <= 12'h603;
      20'h0cf54: out <= 12'h603;
      20'h0cf55: out <= 12'h603;
      20'h0cf56: out <= 12'h603;
      20'h0cf57: out <= 12'h603;
      20'h0cf58: out <= 12'h603;
      20'h0cf59: out <= 12'h603;
      20'h0cf5a: out <= 12'h603;
      20'h0cf5b: out <= 12'h603;
      20'h0cf5c: out <= 12'h603;
      20'h0cf5d: out <= 12'h603;
      20'h0cf5e: out <= 12'h603;
      20'h0cf5f: out <= 12'h603;
      20'h0cf60: out <= 12'h603;
      20'h0cf61: out <= 12'h603;
      20'h0cf62: out <= 12'h603;
      20'h0cf63: out <= 12'h603;
      20'h0cf64: out <= 12'h603;
      20'h0cf65: out <= 12'h603;
      20'h0cf66: out <= 12'h603;
      20'h0cf67: out <= 12'h603;
      20'h0cf68: out <= 12'h603;
      20'h0cf69: out <= 12'h603;
      20'h0cf6a: out <= 12'h603;
      20'h0cf6b: out <= 12'h603;
      20'h0cf6c: out <= 12'h603;
      20'h0cf6d: out <= 12'h603;
      20'h0cf6e: out <= 12'h603;
      20'h0cf6f: out <= 12'h603;
      20'h0cf70: out <= 12'h603;
      20'h0cf71: out <= 12'h603;
      20'h0cf72: out <= 12'h603;
      20'h0cf73: out <= 12'h603;
      20'h0cf74: out <= 12'h603;
      20'h0cf75: out <= 12'h603;
      20'h0cf76: out <= 12'h603;
      20'h0cf77: out <= 12'h603;
      20'h0cf78: out <= 12'h603;
      20'h0cf79: out <= 12'h603;
      20'h0cf7a: out <= 12'h603;
      20'h0cf7b: out <= 12'h603;
      20'h0cf7c: out <= 12'h603;
      20'h0cf7d: out <= 12'h603;
      20'h0cf7e: out <= 12'h603;
      20'h0cf7f: out <= 12'h603;
      20'h0cf80: out <= 12'h603;
      20'h0cf81: out <= 12'h603;
      20'h0cf82: out <= 12'h603;
      20'h0cf83: out <= 12'h603;
      20'h0cf84: out <= 12'h603;
      20'h0cf85: out <= 12'h603;
      20'h0cf86: out <= 12'h603;
      20'h0cf87: out <= 12'h603;
      20'h0cf88: out <= 12'h603;
      20'h0cf89: out <= 12'h603;
      20'h0cf8a: out <= 12'h603;
      20'h0cf8b: out <= 12'h603;
      20'h0cf8c: out <= 12'h603;
      20'h0cf8d: out <= 12'h603;
      20'h0cf8e: out <= 12'h603;
      20'h0cf8f: out <= 12'h603;
      20'h0cf90: out <= 12'hee9;
      20'h0cf91: out <= 12'hf87;
      20'h0cf92: out <= 12'hee9;
      20'h0cf93: out <= 12'hb27;
      20'h0cf94: out <= 12'hb27;
      20'h0cf95: out <= 12'hb27;
      20'h0cf96: out <= 12'hf87;
      20'h0cf97: out <= 12'hb27;
      20'h0cf98: out <= 12'h000;
      20'h0cf99: out <= 12'h000;
      20'h0cf9a: out <= 12'h000;
      20'h0cf9b: out <= 12'h000;
      20'h0cf9c: out <= 12'h000;
      20'h0cf9d: out <= 12'h000;
      20'h0cf9e: out <= 12'h000;
      20'h0cf9f: out <= 12'h000;
      20'h0cfa0: out <= 12'h000;
      20'h0cfa1: out <= 12'h000;
      20'h0cfa2: out <= 12'h000;
      20'h0cfa3: out <= 12'h000;
      20'h0cfa4: out <= 12'h000;
      20'h0cfa5: out <= 12'h000;
      20'h0cfa6: out <= 12'h000;
      20'h0cfa7: out <= 12'h000;
      20'h0cfa8: out <= 12'h000;
      20'h0cfa9: out <= 12'h000;
      20'h0cfaa: out <= 12'h000;
      20'h0cfab: out <= 12'h000;
      20'h0cfac: out <= 12'h000;
      20'h0cfad: out <= 12'h000;
      20'h0cfae: out <= 12'h000;
      20'h0cfaf: out <= 12'h000;
      20'h0cfb0: out <= 12'h000;
      20'h0cfb1: out <= 12'h000;
      20'h0cfb2: out <= 12'h000;
      20'h0cfb3: out <= 12'h000;
      20'h0cfb4: out <= 12'h000;
      20'h0cfb5: out <= 12'h000;
      20'h0cfb6: out <= 12'h000;
      20'h0cfb7: out <= 12'h000;
      20'h0cfb8: out <= 12'h000;
      20'h0cfb9: out <= 12'h000;
      20'h0cfba: out <= 12'h000;
      20'h0cfbb: out <= 12'h000;
      20'h0cfbc: out <= 12'h000;
      20'h0cfbd: out <= 12'h000;
      20'h0cfbe: out <= 12'h000;
      20'h0cfbf: out <= 12'h000;
      20'h0cfc0: out <= 12'h000;
      20'h0cfc1: out <= 12'h000;
      20'h0cfc2: out <= 12'h000;
      20'h0cfc3: out <= 12'h000;
      20'h0cfc4: out <= 12'h000;
      20'h0cfc5: out <= 12'h000;
      20'h0cfc6: out <= 12'h000;
      20'h0cfc7: out <= 12'h000;
      20'h0cfc8: out <= 12'h000;
      20'h0cfc9: out <= 12'h000;
      20'h0cfca: out <= 12'h000;
      20'h0cfcb: out <= 12'h000;
      20'h0cfcc: out <= 12'h000;
      20'h0cfcd: out <= 12'h000;
      20'h0cfce: out <= 12'h000;
      20'h0cfcf: out <= 12'h000;
      20'h0cfd0: out <= 12'h088;
      20'h0cfd1: out <= 12'h088;
      20'h0cfd2: out <= 12'h088;
      20'h0cfd3: out <= 12'h088;
      20'h0cfd4: out <= 12'h088;
      20'h0cfd5: out <= 12'h088;
      20'h0cfd6: out <= 12'h088;
      20'h0cfd7: out <= 12'h088;
      20'h0cfd8: out <= 12'h088;
      20'h0cfd9: out <= 12'h088;
      20'h0cfda: out <= 12'h088;
      20'h0cfdb: out <= 12'h088;
      20'h0cfdc: out <= 12'h088;
      20'h0cfdd: out <= 12'h088;
      20'h0cfde: out <= 12'h088;
      20'h0cfdf: out <= 12'h088;
      20'h0cfe0: out <= 12'h088;
      20'h0cfe1: out <= 12'h088;
      20'h0cfe2: out <= 12'h088;
      20'h0cfe3: out <= 12'h088;
      20'h0cfe4: out <= 12'h088;
      20'h0cfe5: out <= 12'h088;
      20'h0cfe6: out <= 12'h088;
      20'h0cfe7: out <= 12'h088;
      20'h0cfe8: out <= 12'h088;
      20'h0cfe9: out <= 12'h088;
      20'h0cfea: out <= 12'h088;
      20'h0cfeb: out <= 12'h088;
      20'h0cfec: out <= 12'h088;
      20'h0cfed: out <= 12'h088;
      20'h0cfee: out <= 12'h088;
      20'h0cfef: out <= 12'h088;
      20'h0cff0: out <= 12'h088;
      20'h0cff1: out <= 12'h088;
      20'h0cff2: out <= 12'h088;
      20'h0cff3: out <= 12'h088;
      20'h0cff4: out <= 12'h088;
      20'h0cff5: out <= 12'h088;
      20'h0cff6: out <= 12'h088;
      20'h0cff7: out <= 12'h088;
      20'h0cff8: out <= 12'h088;
      20'h0cff9: out <= 12'h088;
      20'h0cffa: out <= 12'h088;
      20'h0cffb: out <= 12'h088;
      20'h0cffc: out <= 12'h088;
      20'h0cffd: out <= 12'h088;
      20'h0cffe: out <= 12'h088;
      20'h0cfff: out <= 12'h088;
      20'h0d000: out <= 12'h088;
      20'h0d001: out <= 12'h088;
      20'h0d002: out <= 12'h088;
      20'h0d003: out <= 12'h088;
      20'h0d004: out <= 12'h088;
      20'h0d005: out <= 12'h088;
      20'h0d006: out <= 12'h088;
      20'h0d007: out <= 12'h088;
      20'h0d008: out <= 12'h088;
      20'h0d009: out <= 12'h088;
      20'h0d00a: out <= 12'h088;
      20'h0d00b: out <= 12'h088;
      20'h0d00c: out <= 12'h088;
      20'h0d00d: out <= 12'h088;
      20'h0d00e: out <= 12'h088;
      20'h0d00f: out <= 12'h088;
      20'h0d010: out <= 12'h088;
      20'h0d011: out <= 12'h088;
      20'h0d012: out <= 12'h088;
      20'h0d013: out <= 12'h088;
      20'h0d014: out <= 12'h088;
      20'h0d015: out <= 12'h088;
      20'h0d016: out <= 12'h088;
      20'h0d017: out <= 12'h088;
      20'h0d018: out <= 12'h088;
      20'h0d019: out <= 12'h088;
      20'h0d01a: out <= 12'h088;
      20'h0d01b: out <= 12'h088;
      20'h0d01c: out <= 12'h088;
      20'h0d01d: out <= 12'h088;
      20'h0d01e: out <= 12'h088;
      20'h0d01f: out <= 12'h088;
      20'h0d020: out <= 12'h088;
      20'h0d021: out <= 12'h088;
      20'h0d022: out <= 12'h088;
      20'h0d023: out <= 12'h088;
      20'h0d024: out <= 12'h088;
      20'h0d025: out <= 12'h088;
      20'h0d026: out <= 12'h088;
      20'h0d027: out <= 12'h088;
      20'h0d028: out <= 12'h088;
      20'h0d029: out <= 12'h088;
      20'h0d02a: out <= 12'h088;
      20'h0d02b: out <= 12'h088;
      20'h0d02c: out <= 12'h088;
      20'h0d02d: out <= 12'h088;
      20'h0d02e: out <= 12'h088;
      20'h0d02f: out <= 12'h088;
      20'h0d030: out <= 12'h088;
      20'h0d031: out <= 12'h088;
      20'h0d032: out <= 12'h088;
      20'h0d033: out <= 12'h088;
      20'h0d034: out <= 12'h088;
      20'h0d035: out <= 12'h088;
      20'h0d036: out <= 12'h088;
      20'h0d037: out <= 12'h088;
      20'h0d038: out <= 12'h088;
      20'h0d039: out <= 12'h603;
      20'h0d03a: out <= 12'h603;
      20'h0d03b: out <= 12'h603;
      20'h0d03c: out <= 12'h603;
      20'h0d03d: out <= 12'h603;
      20'h0d03e: out <= 12'h603;
      20'h0d03f: out <= 12'h603;
      20'h0d040: out <= 12'h603;
      20'h0d041: out <= 12'h603;
      20'h0d042: out <= 12'h603;
      20'h0d043: out <= 12'h603;
      20'h0d044: out <= 12'h603;
      20'h0d045: out <= 12'h603;
      20'h0d046: out <= 12'h603;
      20'h0d047: out <= 12'h603;
      20'h0d048: out <= 12'h603;
      20'h0d049: out <= 12'h603;
      20'h0d04a: out <= 12'h603;
      20'h0d04b: out <= 12'h603;
      20'h0d04c: out <= 12'h603;
      20'h0d04d: out <= 12'h603;
      20'h0d04e: out <= 12'h603;
      20'h0d04f: out <= 12'h603;
      20'h0d050: out <= 12'h603;
      20'h0d051: out <= 12'h603;
      20'h0d052: out <= 12'h603;
      20'h0d053: out <= 12'h603;
      20'h0d054: out <= 12'h603;
      20'h0d055: out <= 12'h603;
      20'h0d056: out <= 12'h603;
      20'h0d057: out <= 12'h603;
      20'h0d058: out <= 12'h603;
      20'h0d059: out <= 12'h603;
      20'h0d05a: out <= 12'h603;
      20'h0d05b: out <= 12'h603;
      20'h0d05c: out <= 12'h603;
      20'h0d05d: out <= 12'h603;
      20'h0d05e: out <= 12'h603;
      20'h0d05f: out <= 12'h603;
      20'h0d060: out <= 12'h603;
      20'h0d061: out <= 12'h603;
      20'h0d062: out <= 12'h603;
      20'h0d063: out <= 12'h603;
      20'h0d064: out <= 12'h603;
      20'h0d065: out <= 12'h603;
      20'h0d066: out <= 12'h603;
      20'h0d067: out <= 12'h603;
      20'h0d068: out <= 12'h603;
      20'h0d069: out <= 12'h603;
      20'h0d06a: out <= 12'h603;
      20'h0d06b: out <= 12'h603;
      20'h0d06c: out <= 12'h603;
      20'h0d06d: out <= 12'h603;
      20'h0d06e: out <= 12'h603;
      20'h0d06f: out <= 12'h603;
      20'h0d070: out <= 12'h603;
      20'h0d071: out <= 12'h603;
      20'h0d072: out <= 12'h603;
      20'h0d073: out <= 12'h603;
      20'h0d074: out <= 12'h603;
      20'h0d075: out <= 12'h603;
      20'h0d076: out <= 12'h603;
      20'h0d077: out <= 12'h603;
      20'h0d078: out <= 12'h603;
      20'h0d079: out <= 12'h603;
      20'h0d07a: out <= 12'h603;
      20'h0d07b: out <= 12'h603;
      20'h0d07c: out <= 12'h603;
      20'h0d07d: out <= 12'h603;
      20'h0d07e: out <= 12'h603;
      20'h0d07f: out <= 12'h603;
      20'h0d080: out <= 12'h603;
      20'h0d081: out <= 12'h603;
      20'h0d082: out <= 12'h603;
      20'h0d083: out <= 12'h603;
      20'h0d084: out <= 12'h603;
      20'h0d085: out <= 12'h603;
      20'h0d086: out <= 12'h603;
      20'h0d087: out <= 12'h603;
      20'h0d088: out <= 12'h603;
      20'h0d089: out <= 12'h603;
      20'h0d08a: out <= 12'h603;
      20'h0d08b: out <= 12'h603;
      20'h0d08c: out <= 12'h603;
      20'h0d08d: out <= 12'h603;
      20'h0d08e: out <= 12'h603;
      20'h0d08f: out <= 12'h603;
      20'h0d090: out <= 12'h603;
      20'h0d091: out <= 12'h603;
      20'h0d092: out <= 12'h603;
      20'h0d093: out <= 12'h603;
      20'h0d094: out <= 12'h603;
      20'h0d095: out <= 12'h603;
      20'h0d096: out <= 12'h603;
      20'h0d097: out <= 12'h603;
      20'h0d098: out <= 12'h603;
      20'h0d099: out <= 12'h603;
      20'h0d09a: out <= 12'h603;
      20'h0d09b: out <= 12'h603;
      20'h0d09c: out <= 12'h603;
      20'h0d09d: out <= 12'h603;
      20'h0d09e: out <= 12'h603;
      20'h0d09f: out <= 12'h603;
      20'h0d0a0: out <= 12'h603;
      20'h0d0a1: out <= 12'h603;
      20'h0d0a2: out <= 12'h603;
      20'h0d0a3: out <= 12'h603;
      20'h0d0a4: out <= 12'h603;
      20'h0d0a5: out <= 12'h603;
      20'h0d0a6: out <= 12'h603;
      20'h0d0a7: out <= 12'h603;
      20'h0d0a8: out <= 12'hee9;
      20'h0d0a9: out <= 12'hf87;
      20'h0d0aa: out <= 12'hf87;
      20'h0d0ab: out <= 12'hf87;
      20'h0d0ac: out <= 12'hf87;
      20'h0d0ad: out <= 12'hf87;
      20'h0d0ae: out <= 12'hf87;
      20'h0d0af: out <= 12'hb27;
      20'h0d0b0: out <= 12'h000;
      20'h0d0b1: out <= 12'h000;
      20'h0d0b2: out <= 12'h000;
      20'h0d0b3: out <= 12'h000;
      20'h0d0b4: out <= 12'h000;
      20'h0d0b5: out <= 12'h000;
      20'h0d0b6: out <= 12'h000;
      20'h0d0b7: out <= 12'h000;
      20'h0d0b8: out <= 12'h000;
      20'h0d0b9: out <= 12'h000;
      20'h0d0ba: out <= 12'h000;
      20'h0d0bb: out <= 12'h000;
      20'h0d0bc: out <= 12'h000;
      20'h0d0bd: out <= 12'h000;
      20'h0d0be: out <= 12'h000;
      20'h0d0bf: out <= 12'h000;
      20'h0d0c0: out <= 12'h000;
      20'h0d0c1: out <= 12'h000;
      20'h0d0c2: out <= 12'h000;
      20'h0d0c3: out <= 12'h000;
      20'h0d0c4: out <= 12'h000;
      20'h0d0c5: out <= 12'h000;
      20'h0d0c6: out <= 12'h000;
      20'h0d0c7: out <= 12'h000;
      20'h0d0c8: out <= 12'h000;
      20'h0d0c9: out <= 12'h000;
      20'h0d0ca: out <= 12'h000;
      20'h0d0cb: out <= 12'h000;
      20'h0d0cc: out <= 12'h000;
      20'h0d0cd: out <= 12'h000;
      20'h0d0ce: out <= 12'h000;
      20'h0d0cf: out <= 12'h000;
      20'h0d0d0: out <= 12'h000;
      20'h0d0d1: out <= 12'h000;
      20'h0d0d2: out <= 12'h000;
      20'h0d0d3: out <= 12'h000;
      20'h0d0d4: out <= 12'h000;
      20'h0d0d5: out <= 12'h000;
      20'h0d0d6: out <= 12'h000;
      20'h0d0d7: out <= 12'h000;
      20'h0d0d8: out <= 12'h000;
      20'h0d0d9: out <= 12'h000;
      20'h0d0da: out <= 12'h000;
      20'h0d0db: out <= 12'h000;
      20'h0d0dc: out <= 12'h000;
      20'h0d0dd: out <= 12'h000;
      20'h0d0de: out <= 12'h000;
      20'h0d0df: out <= 12'h000;
      20'h0d0e0: out <= 12'h000;
      20'h0d0e1: out <= 12'h000;
      20'h0d0e2: out <= 12'h000;
      20'h0d0e3: out <= 12'h000;
      20'h0d0e4: out <= 12'h000;
      20'h0d0e5: out <= 12'h000;
      20'h0d0e6: out <= 12'h000;
      20'h0d0e7: out <= 12'h000;
      20'h0d0e8: out <= 12'h088;
      20'h0d0e9: out <= 12'h088;
      20'h0d0ea: out <= 12'h088;
      20'h0d0eb: out <= 12'h088;
      20'h0d0ec: out <= 12'h088;
      20'h0d0ed: out <= 12'h088;
      20'h0d0ee: out <= 12'h088;
      20'h0d0ef: out <= 12'h088;
      20'h0d0f0: out <= 12'h088;
      20'h0d0f1: out <= 12'h088;
      20'h0d0f2: out <= 12'h088;
      20'h0d0f3: out <= 12'h088;
      20'h0d0f4: out <= 12'h088;
      20'h0d0f5: out <= 12'h088;
      20'h0d0f6: out <= 12'h088;
      20'h0d0f7: out <= 12'h088;
      20'h0d0f8: out <= 12'h088;
      20'h0d0f9: out <= 12'h088;
      20'h0d0fa: out <= 12'h088;
      20'h0d0fb: out <= 12'h088;
      20'h0d0fc: out <= 12'h088;
      20'h0d0fd: out <= 12'h088;
      20'h0d0fe: out <= 12'h088;
      20'h0d0ff: out <= 12'h088;
      20'h0d100: out <= 12'h088;
      20'h0d101: out <= 12'h088;
      20'h0d102: out <= 12'h088;
      20'h0d103: out <= 12'h088;
      20'h0d104: out <= 12'h088;
      20'h0d105: out <= 12'h088;
      20'h0d106: out <= 12'h088;
      20'h0d107: out <= 12'h088;
      20'h0d108: out <= 12'h088;
      20'h0d109: out <= 12'h088;
      20'h0d10a: out <= 12'h088;
      20'h0d10b: out <= 12'h088;
      20'h0d10c: out <= 12'h088;
      20'h0d10d: out <= 12'h088;
      20'h0d10e: out <= 12'h088;
      20'h0d10f: out <= 12'h088;
      20'h0d110: out <= 12'h088;
      20'h0d111: out <= 12'h088;
      20'h0d112: out <= 12'h088;
      20'h0d113: out <= 12'h088;
      20'h0d114: out <= 12'h088;
      20'h0d115: out <= 12'h088;
      20'h0d116: out <= 12'h088;
      20'h0d117: out <= 12'h088;
      20'h0d118: out <= 12'h088;
      20'h0d119: out <= 12'h088;
      20'h0d11a: out <= 12'h088;
      20'h0d11b: out <= 12'h088;
      20'h0d11c: out <= 12'h088;
      20'h0d11d: out <= 12'h088;
      20'h0d11e: out <= 12'h088;
      20'h0d11f: out <= 12'h088;
      20'h0d120: out <= 12'h088;
      20'h0d121: out <= 12'h088;
      20'h0d122: out <= 12'h088;
      20'h0d123: out <= 12'h088;
      20'h0d124: out <= 12'h088;
      20'h0d125: out <= 12'h088;
      20'h0d126: out <= 12'h088;
      20'h0d127: out <= 12'h088;
      20'h0d128: out <= 12'h088;
      20'h0d129: out <= 12'h088;
      20'h0d12a: out <= 12'h088;
      20'h0d12b: out <= 12'h088;
      20'h0d12c: out <= 12'h088;
      20'h0d12d: out <= 12'h088;
      20'h0d12e: out <= 12'h088;
      20'h0d12f: out <= 12'h088;
      20'h0d130: out <= 12'h088;
      20'h0d131: out <= 12'h088;
      20'h0d132: out <= 12'h088;
      20'h0d133: out <= 12'h088;
      20'h0d134: out <= 12'h088;
      20'h0d135: out <= 12'h088;
      20'h0d136: out <= 12'h088;
      20'h0d137: out <= 12'h088;
      20'h0d138: out <= 12'h088;
      20'h0d139: out <= 12'h088;
      20'h0d13a: out <= 12'h088;
      20'h0d13b: out <= 12'h088;
      20'h0d13c: out <= 12'h088;
      20'h0d13d: out <= 12'h088;
      20'h0d13e: out <= 12'h088;
      20'h0d13f: out <= 12'h088;
      20'h0d140: out <= 12'h088;
      20'h0d141: out <= 12'h088;
      20'h0d142: out <= 12'h088;
      20'h0d143: out <= 12'h088;
      20'h0d144: out <= 12'h088;
      20'h0d145: out <= 12'h088;
      20'h0d146: out <= 12'h088;
      20'h0d147: out <= 12'h088;
      20'h0d148: out <= 12'h088;
      20'h0d149: out <= 12'h088;
      20'h0d14a: out <= 12'h088;
      20'h0d14b: out <= 12'h088;
      20'h0d14c: out <= 12'h088;
      20'h0d14d: out <= 12'h088;
      20'h0d14e: out <= 12'h088;
      20'h0d14f: out <= 12'h088;
      20'h0d150: out <= 12'h088;
      20'h0d151: out <= 12'h603;
      20'h0d152: out <= 12'h603;
      20'h0d153: out <= 12'h603;
      20'h0d154: out <= 12'h603;
      20'h0d155: out <= 12'h603;
      20'h0d156: out <= 12'h603;
      20'h0d157: out <= 12'h603;
      20'h0d158: out <= 12'h603;
      20'h0d159: out <= 12'h603;
      20'h0d15a: out <= 12'h603;
      20'h0d15b: out <= 12'h603;
      20'h0d15c: out <= 12'h603;
      20'h0d15d: out <= 12'h603;
      20'h0d15e: out <= 12'h603;
      20'h0d15f: out <= 12'h603;
      20'h0d160: out <= 12'h603;
      20'h0d161: out <= 12'h603;
      20'h0d162: out <= 12'h603;
      20'h0d163: out <= 12'h603;
      20'h0d164: out <= 12'h603;
      20'h0d165: out <= 12'h603;
      20'h0d166: out <= 12'h603;
      20'h0d167: out <= 12'h603;
      20'h0d168: out <= 12'h603;
      20'h0d169: out <= 12'h603;
      20'h0d16a: out <= 12'h603;
      20'h0d16b: out <= 12'h603;
      20'h0d16c: out <= 12'h603;
      20'h0d16d: out <= 12'h603;
      20'h0d16e: out <= 12'h603;
      20'h0d16f: out <= 12'h603;
      20'h0d170: out <= 12'h603;
      20'h0d171: out <= 12'h603;
      20'h0d172: out <= 12'h603;
      20'h0d173: out <= 12'h603;
      20'h0d174: out <= 12'h603;
      20'h0d175: out <= 12'h603;
      20'h0d176: out <= 12'h603;
      20'h0d177: out <= 12'h603;
      20'h0d178: out <= 12'h603;
      20'h0d179: out <= 12'h603;
      20'h0d17a: out <= 12'h603;
      20'h0d17b: out <= 12'h603;
      20'h0d17c: out <= 12'h603;
      20'h0d17d: out <= 12'h603;
      20'h0d17e: out <= 12'h603;
      20'h0d17f: out <= 12'h603;
      20'h0d180: out <= 12'h603;
      20'h0d181: out <= 12'h603;
      20'h0d182: out <= 12'h603;
      20'h0d183: out <= 12'h603;
      20'h0d184: out <= 12'h603;
      20'h0d185: out <= 12'h603;
      20'h0d186: out <= 12'h603;
      20'h0d187: out <= 12'h603;
      20'h0d188: out <= 12'h603;
      20'h0d189: out <= 12'h603;
      20'h0d18a: out <= 12'h603;
      20'h0d18b: out <= 12'h603;
      20'h0d18c: out <= 12'h603;
      20'h0d18d: out <= 12'h603;
      20'h0d18e: out <= 12'h603;
      20'h0d18f: out <= 12'h603;
      20'h0d190: out <= 12'h603;
      20'h0d191: out <= 12'h603;
      20'h0d192: out <= 12'h603;
      20'h0d193: out <= 12'h603;
      20'h0d194: out <= 12'h603;
      20'h0d195: out <= 12'h603;
      20'h0d196: out <= 12'h603;
      20'h0d197: out <= 12'h603;
      20'h0d198: out <= 12'h603;
      20'h0d199: out <= 12'h603;
      20'h0d19a: out <= 12'h603;
      20'h0d19b: out <= 12'h603;
      20'h0d19c: out <= 12'h603;
      20'h0d19d: out <= 12'h603;
      20'h0d19e: out <= 12'h603;
      20'h0d19f: out <= 12'h603;
      20'h0d1a0: out <= 12'h603;
      20'h0d1a1: out <= 12'h603;
      20'h0d1a2: out <= 12'h603;
      20'h0d1a3: out <= 12'h603;
      20'h0d1a4: out <= 12'h603;
      20'h0d1a5: out <= 12'h603;
      20'h0d1a6: out <= 12'h603;
      20'h0d1a7: out <= 12'h603;
      20'h0d1a8: out <= 12'h603;
      20'h0d1a9: out <= 12'h603;
      20'h0d1aa: out <= 12'h603;
      20'h0d1ab: out <= 12'h603;
      20'h0d1ac: out <= 12'h603;
      20'h0d1ad: out <= 12'h603;
      20'h0d1ae: out <= 12'h603;
      20'h0d1af: out <= 12'h603;
      20'h0d1b0: out <= 12'h603;
      20'h0d1b1: out <= 12'h603;
      20'h0d1b2: out <= 12'h603;
      20'h0d1b3: out <= 12'h603;
      20'h0d1b4: out <= 12'h603;
      20'h0d1b5: out <= 12'h603;
      20'h0d1b6: out <= 12'h603;
      20'h0d1b7: out <= 12'h603;
      20'h0d1b8: out <= 12'h603;
      20'h0d1b9: out <= 12'h603;
      20'h0d1ba: out <= 12'h603;
      20'h0d1bb: out <= 12'h603;
      20'h0d1bc: out <= 12'h603;
      20'h0d1bd: out <= 12'h603;
      20'h0d1be: out <= 12'h603;
      20'h0d1bf: out <= 12'h603;
      20'h0d1c0: out <= 12'hb27;
      20'h0d1c1: out <= 12'hb27;
      20'h0d1c2: out <= 12'hb27;
      20'h0d1c3: out <= 12'hb27;
      20'h0d1c4: out <= 12'hb27;
      20'h0d1c5: out <= 12'hb27;
      20'h0d1c6: out <= 12'hb27;
      20'h0d1c7: out <= 12'hb27;
      20'h0d1c8: out <= 12'h000;
      20'h0d1c9: out <= 12'h000;
      20'h0d1ca: out <= 12'h000;
      20'h0d1cb: out <= 12'h000;
      20'h0d1cc: out <= 12'h000;
      20'h0d1cd: out <= 12'h000;
      20'h0d1ce: out <= 12'h000;
      20'h0d1cf: out <= 12'h000;
      20'h0d1d0: out <= 12'h000;
      20'h0d1d1: out <= 12'h000;
      20'h0d1d2: out <= 12'h000;
      20'h0d1d3: out <= 12'h000;
      20'h0d1d4: out <= 12'h000;
      20'h0d1d5: out <= 12'h000;
      20'h0d1d6: out <= 12'h000;
      20'h0d1d7: out <= 12'h000;
      20'h0d1d8: out <= 12'h000;
      20'h0d1d9: out <= 12'h000;
      20'h0d1da: out <= 12'h000;
      20'h0d1db: out <= 12'h000;
      20'h0d1dc: out <= 12'h000;
      20'h0d1dd: out <= 12'h000;
      20'h0d1de: out <= 12'h000;
      20'h0d1df: out <= 12'h000;
      20'h0d1e0: out <= 12'h000;
      20'h0d1e1: out <= 12'h000;
      20'h0d1e2: out <= 12'h000;
      20'h0d1e3: out <= 12'h000;
      20'h0d1e4: out <= 12'h000;
      20'h0d1e5: out <= 12'h000;
      20'h0d1e6: out <= 12'h000;
      20'h0d1e7: out <= 12'h000;
      20'h0d1e8: out <= 12'h000;
      20'h0d1e9: out <= 12'h000;
      20'h0d1ea: out <= 12'h000;
      20'h0d1eb: out <= 12'h000;
      20'h0d1ec: out <= 12'h000;
      20'h0d1ed: out <= 12'h000;
      20'h0d1ee: out <= 12'h000;
      20'h0d1ef: out <= 12'h000;
      20'h0d1f0: out <= 12'h000;
      20'h0d1f1: out <= 12'h000;
      20'h0d1f2: out <= 12'h000;
      20'h0d1f3: out <= 12'h000;
      20'h0d1f4: out <= 12'h000;
      20'h0d1f5: out <= 12'h000;
      20'h0d1f6: out <= 12'h000;
      20'h0d1f7: out <= 12'h000;
      20'h0d1f8: out <= 12'h000;
      20'h0d1f9: out <= 12'h000;
      20'h0d1fa: out <= 12'h000;
      20'h0d1fb: out <= 12'h000;
      20'h0d1fc: out <= 12'h000;
      20'h0d1fd: out <= 12'h000;
      20'h0d1fe: out <= 12'h000;
      20'h0d1ff: out <= 12'h000;
      20'h0d200: out <= 12'h088;
      20'h0d201: out <= 12'h088;
      20'h0d202: out <= 12'h088;
      20'h0d203: out <= 12'h088;
      20'h0d204: out <= 12'h088;
      20'h0d205: out <= 12'h088;
      20'h0d206: out <= 12'h088;
      20'h0d207: out <= 12'h088;
      20'h0d208: out <= 12'h088;
      20'h0d209: out <= 12'h088;
      20'h0d20a: out <= 12'h088;
      20'h0d20b: out <= 12'h088;
      20'h0d20c: out <= 12'h088;
      20'h0d20d: out <= 12'h088;
      20'h0d20e: out <= 12'h088;
      20'h0d20f: out <= 12'h088;
      20'h0d210: out <= 12'h088;
      20'h0d211: out <= 12'h088;
      20'h0d212: out <= 12'h088;
      20'h0d213: out <= 12'h088;
      20'h0d214: out <= 12'h088;
      20'h0d215: out <= 12'h088;
      20'h0d216: out <= 12'h088;
      20'h0d217: out <= 12'h088;
      20'h0d218: out <= 12'h088;
      20'h0d219: out <= 12'h088;
      20'h0d21a: out <= 12'h088;
      20'h0d21b: out <= 12'h088;
      20'h0d21c: out <= 12'h088;
      20'h0d21d: out <= 12'h088;
      20'h0d21e: out <= 12'h088;
      20'h0d21f: out <= 12'h088;
      20'h0d220: out <= 12'h088;
      20'h0d221: out <= 12'h088;
      20'h0d222: out <= 12'h088;
      20'h0d223: out <= 12'h088;
      20'h0d224: out <= 12'h088;
      20'h0d225: out <= 12'h088;
      20'h0d226: out <= 12'h088;
      20'h0d227: out <= 12'h088;
      20'h0d228: out <= 12'h088;
      20'h0d229: out <= 12'h088;
      20'h0d22a: out <= 12'h088;
      20'h0d22b: out <= 12'h088;
      20'h0d22c: out <= 12'h088;
      20'h0d22d: out <= 12'h088;
      20'h0d22e: out <= 12'h088;
      20'h0d22f: out <= 12'h088;
      20'h0d230: out <= 12'h088;
      20'h0d231: out <= 12'h088;
      20'h0d232: out <= 12'h088;
      20'h0d233: out <= 12'h088;
      20'h0d234: out <= 12'h088;
      20'h0d235: out <= 12'h088;
      20'h0d236: out <= 12'h088;
      20'h0d237: out <= 12'h088;
      20'h0d238: out <= 12'h088;
      20'h0d239: out <= 12'h088;
      20'h0d23a: out <= 12'h088;
      20'h0d23b: out <= 12'h088;
      20'h0d23c: out <= 12'h088;
      20'h0d23d: out <= 12'h088;
      20'h0d23e: out <= 12'h088;
      20'h0d23f: out <= 12'h088;
      20'h0d240: out <= 12'h088;
      20'h0d241: out <= 12'h088;
      20'h0d242: out <= 12'h088;
      20'h0d243: out <= 12'h088;
      20'h0d244: out <= 12'h088;
      20'h0d245: out <= 12'h088;
      20'h0d246: out <= 12'h088;
      20'h0d247: out <= 12'h088;
      20'h0d248: out <= 12'h088;
      20'h0d249: out <= 12'h088;
      20'h0d24a: out <= 12'h088;
      20'h0d24b: out <= 12'h088;
      20'h0d24c: out <= 12'h088;
      20'h0d24d: out <= 12'h088;
      20'h0d24e: out <= 12'h088;
      20'h0d24f: out <= 12'h088;
      20'h0d250: out <= 12'h088;
      20'h0d251: out <= 12'h088;
      20'h0d252: out <= 12'h088;
      20'h0d253: out <= 12'h088;
      20'h0d254: out <= 12'h088;
      20'h0d255: out <= 12'h088;
      20'h0d256: out <= 12'h088;
      20'h0d257: out <= 12'h088;
      20'h0d258: out <= 12'h088;
      20'h0d259: out <= 12'h088;
      20'h0d25a: out <= 12'h088;
      20'h0d25b: out <= 12'h088;
      20'h0d25c: out <= 12'h088;
      20'h0d25d: out <= 12'h088;
      20'h0d25e: out <= 12'h088;
      20'h0d25f: out <= 12'h088;
      20'h0d260: out <= 12'h088;
      20'h0d261: out <= 12'h088;
      20'h0d262: out <= 12'h088;
      20'h0d263: out <= 12'h088;
      20'h0d264: out <= 12'h088;
      20'h0d265: out <= 12'h088;
      20'h0d266: out <= 12'h088;
      20'h0d267: out <= 12'h088;
      20'h0d268: out <= 12'h088;
      20'h0d269: out <= 12'h000;
      20'h0d26a: out <= 12'h000;
      20'h0d26b: out <= 12'h000;
      20'h0d26c: out <= 12'h000;
      20'h0d26d: out <= 12'h000;
      20'h0d26e: out <= 12'h000;
      20'h0d26f: out <= 12'h000;
      20'h0d270: out <= 12'h000;
      20'h0d271: out <= 12'h000;
      20'h0d272: out <= 12'h000;
      20'h0d273: out <= 12'h000;
      20'h0d274: out <= 12'h000;
      20'h0d275: out <= 12'h000;
      20'h0d276: out <= 12'h000;
      20'h0d277: out <= 12'h000;
      20'h0d278: out <= 12'h000;
      20'h0d279: out <= 12'h000;
      20'h0d27a: out <= 12'h000;
      20'h0d27b: out <= 12'h000;
      20'h0d27c: out <= 12'h000;
      20'h0d27d: out <= 12'h000;
      20'h0d27e: out <= 12'h000;
      20'h0d27f: out <= 12'h000;
      20'h0d280: out <= 12'h603;
      20'h0d281: out <= 12'h603;
      20'h0d282: out <= 12'h603;
      20'h0d283: out <= 12'h603;
      20'h0d284: out <= 12'h603;
      20'h0d285: out <= 12'h603;
      20'h0d286: out <= 12'h603;
      20'h0d287: out <= 12'h603;
      20'h0d288: out <= 12'h603;
      20'h0d289: out <= 12'h603;
      20'h0d28a: out <= 12'h603;
      20'h0d28b: out <= 12'h603;
      20'h0d28c: out <= 12'h603;
      20'h0d28d: out <= 12'h603;
      20'h0d28e: out <= 12'h603;
      20'h0d28f: out <= 12'h603;
      20'h0d290: out <= 12'h603;
      20'h0d291: out <= 12'h603;
      20'h0d292: out <= 12'h603;
      20'h0d293: out <= 12'h603;
      20'h0d294: out <= 12'h603;
      20'h0d295: out <= 12'h603;
      20'h0d296: out <= 12'h603;
      20'h0d297: out <= 12'h603;
      20'h0d298: out <= 12'h603;
      20'h0d299: out <= 12'h603;
      20'h0d29a: out <= 12'h603;
      20'h0d29b: out <= 12'h603;
      20'h0d29c: out <= 12'h603;
      20'h0d29d: out <= 12'h603;
      20'h0d29e: out <= 12'h603;
      20'h0d29f: out <= 12'h603;
      20'h0d2a0: out <= 12'h603;
      20'h0d2a1: out <= 12'h603;
      20'h0d2a2: out <= 12'h603;
      20'h0d2a3: out <= 12'h603;
      20'h0d2a4: out <= 12'h603;
      20'h0d2a5: out <= 12'h603;
      20'h0d2a6: out <= 12'h603;
      20'h0d2a7: out <= 12'h603;
      20'h0d2a8: out <= 12'h603;
      20'h0d2a9: out <= 12'h603;
      20'h0d2aa: out <= 12'h603;
      20'h0d2ab: out <= 12'h603;
      20'h0d2ac: out <= 12'h603;
      20'h0d2ad: out <= 12'h603;
      20'h0d2ae: out <= 12'h603;
      20'h0d2af: out <= 12'h603;
      20'h0d2b0: out <= 12'h603;
      20'h0d2b1: out <= 12'h603;
      20'h0d2b2: out <= 12'h603;
      20'h0d2b3: out <= 12'h603;
      20'h0d2b4: out <= 12'h603;
      20'h0d2b5: out <= 12'h603;
      20'h0d2b6: out <= 12'h603;
      20'h0d2b7: out <= 12'h603;
      20'h0d2b8: out <= 12'h603;
      20'h0d2b9: out <= 12'h603;
      20'h0d2ba: out <= 12'h603;
      20'h0d2bb: out <= 12'h603;
      20'h0d2bc: out <= 12'h603;
      20'h0d2bd: out <= 12'h603;
      20'h0d2be: out <= 12'h603;
      20'h0d2bf: out <= 12'h603;
      20'h0d2c0: out <= 12'h603;
      20'h0d2c1: out <= 12'h603;
      20'h0d2c2: out <= 12'h603;
      20'h0d2c3: out <= 12'h603;
      20'h0d2c4: out <= 12'h603;
      20'h0d2c5: out <= 12'h603;
      20'h0d2c6: out <= 12'h603;
      20'h0d2c7: out <= 12'h603;
      20'h0d2c8: out <= 12'h603;
      20'h0d2c9: out <= 12'h603;
      20'h0d2ca: out <= 12'h603;
      20'h0d2cb: out <= 12'h603;
      20'h0d2cc: out <= 12'h603;
      20'h0d2cd: out <= 12'h603;
      20'h0d2ce: out <= 12'h603;
      20'h0d2cf: out <= 12'h603;
      20'h0d2d0: out <= 12'h603;
      20'h0d2d1: out <= 12'h603;
      20'h0d2d2: out <= 12'h603;
      20'h0d2d3: out <= 12'h603;
      20'h0d2d4: out <= 12'h603;
      20'h0d2d5: out <= 12'h603;
      20'h0d2d6: out <= 12'h603;
      20'h0d2d7: out <= 12'h603;
      20'h0d2d8: out <= 12'hee9;
      20'h0d2d9: out <= 12'hee9;
      20'h0d2da: out <= 12'hee9;
      20'h0d2db: out <= 12'hee9;
      20'h0d2dc: out <= 12'hee9;
      20'h0d2dd: out <= 12'hee9;
      20'h0d2de: out <= 12'hee9;
      20'h0d2df: out <= 12'hb27;
      20'h0d2e0: out <= 12'h000;
      20'h0d2e1: out <= 12'h000;
      20'h0d2e2: out <= 12'h000;
      20'h0d2e3: out <= 12'h000;
      20'h0d2e4: out <= 12'h000;
      20'h0d2e5: out <= 12'h000;
      20'h0d2e6: out <= 12'h000;
      20'h0d2e7: out <= 12'h000;
      20'h0d2e8: out <= 12'hbbb;
      20'h0d2e9: out <= 12'hbbb;
      20'h0d2ea: out <= 12'hbbb;
      20'h0d2eb: out <= 12'hbbb;
      20'h0d2ec: out <= 12'hbbb;
      20'h0d2ed: out <= 12'h000;
      20'h0d2ee: out <= 12'h000;
      20'h0d2ef: out <= 12'hbbb;
      20'h0d2f0: out <= 12'hbbb;
      20'h0d2f1: out <= 12'hbbb;
      20'h0d2f2: out <= 12'hbbb;
      20'h0d2f3: out <= 12'h000;
      20'h0d2f4: out <= 12'h000;
      20'h0d2f5: out <= 12'hbbb;
      20'h0d2f6: out <= 12'hbbb;
      20'h0d2f7: out <= 12'hbbb;
      20'h0d2f8: out <= 12'hbbb;
      20'h0d2f9: out <= 12'hbbb;
      20'h0d2fa: out <= 12'h000;
      20'h0d2fb: out <= 12'h000;
      20'h0d2fc: out <= 12'hbbb;
      20'h0d2fd: out <= 12'hbbb;
      20'h0d2fe: out <= 12'hbbb;
      20'h0d2ff: out <= 12'h000;
      20'h0d300: out <= 12'hbbb;
      20'h0d301: out <= 12'hbbb;
      20'h0d302: out <= 12'h000;
      20'h0d303: out <= 12'h000;
      20'h0d304: out <= 12'hbbb;
      20'h0d305: out <= 12'hbbb;
      20'h0d306: out <= 12'h000;
      20'h0d307: out <= 12'h000;
      20'h0d308: out <= 12'h000;
      20'h0d309: out <= 12'hbbb;
      20'h0d30a: out <= 12'hbbb;
      20'h0d30b: out <= 12'h000;
      20'h0d30c: out <= 12'h000;
      20'h0d30d: out <= 12'h000;
      20'h0d30e: out <= 12'h000;
      20'h0d30f: out <= 12'h000;
      20'h0d310: out <= 12'h000;
      20'h0d311: out <= 12'h000;
      20'h0d312: out <= 12'h000;
      20'h0d313: out <= 12'h000;
      20'h0d314: out <= 12'h000;
      20'h0d315: out <= 12'h000;
      20'h0d316: out <= 12'h000;
      20'h0d317: out <= 12'h000;
      20'h0d318: out <= 12'h088;
      20'h0d319: out <= 12'h088;
      20'h0d31a: out <= 12'h088;
      20'h0d31b: out <= 12'h088;
      20'h0d31c: out <= 12'h088;
      20'h0d31d: out <= 12'h088;
      20'h0d31e: out <= 12'h088;
      20'h0d31f: out <= 12'h088;
      20'h0d320: out <= 12'h088;
      20'h0d321: out <= 12'h088;
      20'h0d322: out <= 12'h088;
      20'h0d323: out <= 12'h088;
      20'h0d324: out <= 12'h088;
      20'h0d325: out <= 12'h088;
      20'h0d326: out <= 12'h088;
      20'h0d327: out <= 12'h088;
      20'h0d328: out <= 12'h088;
      20'h0d329: out <= 12'h088;
      20'h0d32a: out <= 12'h088;
      20'h0d32b: out <= 12'h088;
      20'h0d32c: out <= 12'h088;
      20'h0d32d: out <= 12'h088;
      20'h0d32e: out <= 12'h088;
      20'h0d32f: out <= 12'h088;
      20'h0d330: out <= 12'h088;
      20'h0d331: out <= 12'h088;
      20'h0d332: out <= 12'h088;
      20'h0d333: out <= 12'h088;
      20'h0d334: out <= 12'h088;
      20'h0d335: out <= 12'h088;
      20'h0d336: out <= 12'h088;
      20'h0d337: out <= 12'h088;
      20'h0d338: out <= 12'h088;
      20'h0d339: out <= 12'h088;
      20'h0d33a: out <= 12'h088;
      20'h0d33b: out <= 12'h088;
      20'h0d33c: out <= 12'h088;
      20'h0d33d: out <= 12'h088;
      20'h0d33e: out <= 12'h088;
      20'h0d33f: out <= 12'h088;
      20'h0d340: out <= 12'h088;
      20'h0d341: out <= 12'h088;
      20'h0d342: out <= 12'h088;
      20'h0d343: out <= 12'h088;
      20'h0d344: out <= 12'h088;
      20'h0d345: out <= 12'h088;
      20'h0d346: out <= 12'h088;
      20'h0d347: out <= 12'h088;
      20'h0d348: out <= 12'h088;
      20'h0d349: out <= 12'h088;
      20'h0d34a: out <= 12'h088;
      20'h0d34b: out <= 12'h088;
      20'h0d34c: out <= 12'h088;
      20'h0d34d: out <= 12'h088;
      20'h0d34e: out <= 12'h088;
      20'h0d34f: out <= 12'h088;
      20'h0d350: out <= 12'h088;
      20'h0d351: out <= 12'h088;
      20'h0d352: out <= 12'h088;
      20'h0d353: out <= 12'h088;
      20'h0d354: out <= 12'h088;
      20'h0d355: out <= 12'h088;
      20'h0d356: out <= 12'h088;
      20'h0d357: out <= 12'h088;
      20'h0d358: out <= 12'h088;
      20'h0d359: out <= 12'h088;
      20'h0d35a: out <= 12'h088;
      20'h0d35b: out <= 12'h088;
      20'h0d35c: out <= 12'h088;
      20'h0d35d: out <= 12'h088;
      20'h0d35e: out <= 12'h088;
      20'h0d35f: out <= 12'h088;
      20'h0d360: out <= 12'h088;
      20'h0d361: out <= 12'h088;
      20'h0d362: out <= 12'h088;
      20'h0d363: out <= 12'h088;
      20'h0d364: out <= 12'h088;
      20'h0d365: out <= 12'h088;
      20'h0d366: out <= 12'h088;
      20'h0d367: out <= 12'h088;
      20'h0d368: out <= 12'h088;
      20'h0d369: out <= 12'h088;
      20'h0d36a: out <= 12'h088;
      20'h0d36b: out <= 12'h088;
      20'h0d36c: out <= 12'h088;
      20'h0d36d: out <= 12'h088;
      20'h0d36e: out <= 12'h088;
      20'h0d36f: out <= 12'h088;
      20'h0d370: out <= 12'h088;
      20'h0d371: out <= 12'h088;
      20'h0d372: out <= 12'h088;
      20'h0d373: out <= 12'h088;
      20'h0d374: out <= 12'h088;
      20'h0d375: out <= 12'h088;
      20'h0d376: out <= 12'h088;
      20'h0d377: out <= 12'h088;
      20'h0d378: out <= 12'h088;
      20'h0d379: out <= 12'h088;
      20'h0d37a: out <= 12'h088;
      20'h0d37b: out <= 12'h088;
      20'h0d37c: out <= 12'h088;
      20'h0d37d: out <= 12'h088;
      20'h0d37e: out <= 12'h088;
      20'h0d37f: out <= 12'h088;
      20'h0d380: out <= 12'h088;
      20'h0d381: out <= 12'h6af;
      20'h0d382: out <= 12'h6af;
      20'h0d383: out <= 12'h16d;
      20'h0d384: out <= 12'h16d;
      20'h0d385: out <= 12'h16d;
      20'h0d386: out <= 12'h000;
      20'h0d387: out <= 12'h000;
      20'h0d388: out <= 12'h000;
      20'h0d389: out <= 12'h000;
      20'h0d38a: out <= 12'h660;
      20'h0d38b: out <= 12'h660;
      20'h0d38c: out <= 12'h660;
      20'h0d38d: out <= 12'hbb0;
      20'h0d38e: out <= 12'hbb0;
      20'h0d38f: out <= 12'hbb0;
      20'h0d390: out <= 12'hbb0;
      20'h0d391: out <= 12'hbb0;
      20'h0d392: out <= 12'hbb0;
      20'h0d393: out <= 12'h660;
      20'h0d394: out <= 12'h660;
      20'h0d395: out <= 12'h660;
      20'h0d396: out <= 12'h000;
      20'h0d397: out <= 12'h000;
      20'h0d398: out <= 12'h603;
      20'h0d399: out <= 12'h603;
      20'h0d39a: out <= 12'h603;
      20'h0d39b: out <= 12'h603;
      20'h0d39c: out <= 12'h603;
      20'h0d39d: out <= 12'h603;
      20'h0d39e: out <= 12'h603;
      20'h0d39f: out <= 12'h603;
      20'h0d3a0: out <= 12'h603;
      20'h0d3a1: out <= 12'h603;
      20'h0d3a2: out <= 12'h603;
      20'h0d3a3: out <= 12'h603;
      20'h0d3a4: out <= 12'h603;
      20'h0d3a5: out <= 12'h603;
      20'h0d3a6: out <= 12'h603;
      20'h0d3a7: out <= 12'h603;
      20'h0d3a8: out <= 12'h603;
      20'h0d3a9: out <= 12'h603;
      20'h0d3aa: out <= 12'h603;
      20'h0d3ab: out <= 12'h603;
      20'h0d3ac: out <= 12'h603;
      20'h0d3ad: out <= 12'h603;
      20'h0d3ae: out <= 12'h603;
      20'h0d3af: out <= 12'h603;
      20'h0d3b0: out <= 12'h603;
      20'h0d3b1: out <= 12'h603;
      20'h0d3b2: out <= 12'h603;
      20'h0d3b3: out <= 12'h603;
      20'h0d3b4: out <= 12'h603;
      20'h0d3b5: out <= 12'h603;
      20'h0d3b6: out <= 12'h603;
      20'h0d3b7: out <= 12'h603;
      20'h0d3b8: out <= 12'h603;
      20'h0d3b9: out <= 12'h603;
      20'h0d3ba: out <= 12'h603;
      20'h0d3bb: out <= 12'h603;
      20'h0d3bc: out <= 12'h603;
      20'h0d3bd: out <= 12'h603;
      20'h0d3be: out <= 12'h603;
      20'h0d3bf: out <= 12'h603;
      20'h0d3c0: out <= 12'h603;
      20'h0d3c1: out <= 12'h603;
      20'h0d3c2: out <= 12'h603;
      20'h0d3c3: out <= 12'h603;
      20'h0d3c4: out <= 12'h603;
      20'h0d3c5: out <= 12'h603;
      20'h0d3c6: out <= 12'h603;
      20'h0d3c7: out <= 12'h603;
      20'h0d3c8: out <= 12'h603;
      20'h0d3c9: out <= 12'h603;
      20'h0d3ca: out <= 12'h603;
      20'h0d3cb: out <= 12'h603;
      20'h0d3cc: out <= 12'h603;
      20'h0d3cd: out <= 12'h603;
      20'h0d3ce: out <= 12'h603;
      20'h0d3cf: out <= 12'h603;
      20'h0d3d0: out <= 12'h603;
      20'h0d3d1: out <= 12'h603;
      20'h0d3d2: out <= 12'h603;
      20'h0d3d3: out <= 12'h603;
      20'h0d3d4: out <= 12'h603;
      20'h0d3d5: out <= 12'h603;
      20'h0d3d6: out <= 12'h603;
      20'h0d3d7: out <= 12'h603;
      20'h0d3d8: out <= 12'h603;
      20'h0d3d9: out <= 12'h603;
      20'h0d3da: out <= 12'h603;
      20'h0d3db: out <= 12'h603;
      20'h0d3dc: out <= 12'h603;
      20'h0d3dd: out <= 12'h603;
      20'h0d3de: out <= 12'h603;
      20'h0d3df: out <= 12'h603;
      20'h0d3e0: out <= 12'h603;
      20'h0d3e1: out <= 12'h603;
      20'h0d3e2: out <= 12'h603;
      20'h0d3e3: out <= 12'h603;
      20'h0d3e4: out <= 12'h603;
      20'h0d3e5: out <= 12'h603;
      20'h0d3e6: out <= 12'h603;
      20'h0d3e7: out <= 12'h603;
      20'h0d3e8: out <= 12'h603;
      20'h0d3e9: out <= 12'h603;
      20'h0d3ea: out <= 12'h603;
      20'h0d3eb: out <= 12'h603;
      20'h0d3ec: out <= 12'h603;
      20'h0d3ed: out <= 12'h603;
      20'h0d3ee: out <= 12'h603;
      20'h0d3ef: out <= 12'h603;
      20'h0d3f0: out <= 12'hee9;
      20'h0d3f1: out <= 12'hf87;
      20'h0d3f2: out <= 12'hf87;
      20'h0d3f3: out <= 12'hf87;
      20'h0d3f4: out <= 12'hf87;
      20'h0d3f5: out <= 12'hf87;
      20'h0d3f6: out <= 12'hf87;
      20'h0d3f7: out <= 12'hb27;
      20'h0d3f8: out <= 12'h000;
      20'h0d3f9: out <= 12'h000;
      20'h0d3fa: out <= 12'h000;
      20'h0d3fb: out <= 12'h000;
      20'h0d3fc: out <= 12'h000;
      20'h0d3fd: out <= 12'h000;
      20'h0d3fe: out <= 12'h000;
      20'h0d3ff: out <= 12'h000;
      20'h0d400: out <= 12'hbbb;
      20'h0d401: out <= 12'hbbb;
      20'h0d402: out <= 12'h000;
      20'h0d403: out <= 12'h000;
      20'h0d404: out <= 12'h000;
      20'h0d405: out <= 12'h000;
      20'h0d406: out <= 12'hbbb;
      20'h0d407: out <= 12'hbbb;
      20'h0d408: out <= 12'h000;
      20'h0d409: out <= 12'h000;
      20'h0d40a: out <= 12'hbbb;
      20'h0d40b: out <= 12'hbbb;
      20'h0d40c: out <= 12'h000;
      20'h0d40d: out <= 12'hbbb;
      20'h0d40e: out <= 12'hbbb;
      20'h0d40f: out <= 12'h000;
      20'h0d410: out <= 12'h000;
      20'h0d411: out <= 12'h000;
      20'h0d412: out <= 12'h000;
      20'h0d413: out <= 12'hbbb;
      20'h0d414: out <= 12'hbbb;
      20'h0d415: out <= 12'hbbb;
      20'h0d416: out <= 12'hbbb;
      20'h0d417: out <= 12'hbbb;
      20'h0d418: out <= 12'hbbb;
      20'h0d419: out <= 12'hbbb;
      20'h0d41a: out <= 12'hbbb;
      20'h0d41b: out <= 12'h000;
      20'h0d41c: out <= 12'hbbb;
      20'h0d41d: out <= 12'hbbb;
      20'h0d41e: out <= 12'h000;
      20'h0d41f: out <= 12'h000;
      20'h0d420: out <= 12'h000;
      20'h0d421: out <= 12'hbbb;
      20'h0d422: out <= 12'hbbb;
      20'h0d423: out <= 12'h000;
      20'h0d424: out <= 12'h000;
      20'h0d425: out <= 12'h000;
      20'h0d426: out <= 12'h000;
      20'h0d427: out <= 12'h000;
      20'h0d428: out <= 12'h000;
      20'h0d429: out <= 12'h000;
      20'h0d42a: out <= 12'h000;
      20'h0d42b: out <= 12'h000;
      20'h0d42c: out <= 12'h000;
      20'h0d42d: out <= 12'h000;
      20'h0d42e: out <= 12'h000;
      20'h0d42f: out <= 12'h000;
      20'h0d430: out <= 12'h088;
      20'h0d431: out <= 12'h088;
      20'h0d432: out <= 12'h088;
      20'h0d433: out <= 12'h088;
      20'h0d434: out <= 12'h088;
      20'h0d435: out <= 12'h088;
      20'h0d436: out <= 12'h088;
      20'h0d437: out <= 12'h088;
      20'h0d438: out <= 12'h088;
      20'h0d439: out <= 12'h088;
      20'h0d43a: out <= 12'h088;
      20'h0d43b: out <= 12'h088;
      20'h0d43c: out <= 12'h088;
      20'h0d43d: out <= 12'h088;
      20'h0d43e: out <= 12'h088;
      20'h0d43f: out <= 12'h088;
      20'h0d440: out <= 12'h088;
      20'h0d441: out <= 12'h088;
      20'h0d442: out <= 12'h088;
      20'h0d443: out <= 12'h088;
      20'h0d444: out <= 12'h088;
      20'h0d445: out <= 12'h088;
      20'h0d446: out <= 12'h088;
      20'h0d447: out <= 12'h088;
      20'h0d448: out <= 12'h088;
      20'h0d449: out <= 12'h088;
      20'h0d44a: out <= 12'h088;
      20'h0d44b: out <= 12'h088;
      20'h0d44c: out <= 12'h088;
      20'h0d44d: out <= 12'h088;
      20'h0d44e: out <= 12'h088;
      20'h0d44f: out <= 12'h088;
      20'h0d450: out <= 12'h088;
      20'h0d451: out <= 12'h088;
      20'h0d452: out <= 12'h088;
      20'h0d453: out <= 12'h088;
      20'h0d454: out <= 12'h088;
      20'h0d455: out <= 12'h088;
      20'h0d456: out <= 12'h088;
      20'h0d457: out <= 12'h088;
      20'h0d458: out <= 12'h088;
      20'h0d459: out <= 12'h088;
      20'h0d45a: out <= 12'h088;
      20'h0d45b: out <= 12'h088;
      20'h0d45c: out <= 12'h088;
      20'h0d45d: out <= 12'h088;
      20'h0d45e: out <= 12'h088;
      20'h0d45f: out <= 12'h088;
      20'h0d460: out <= 12'h088;
      20'h0d461: out <= 12'h088;
      20'h0d462: out <= 12'h088;
      20'h0d463: out <= 12'h088;
      20'h0d464: out <= 12'h088;
      20'h0d465: out <= 12'h088;
      20'h0d466: out <= 12'h088;
      20'h0d467: out <= 12'h088;
      20'h0d468: out <= 12'h088;
      20'h0d469: out <= 12'h088;
      20'h0d46a: out <= 12'h088;
      20'h0d46b: out <= 12'h088;
      20'h0d46c: out <= 12'h088;
      20'h0d46d: out <= 12'h088;
      20'h0d46e: out <= 12'h088;
      20'h0d46f: out <= 12'h088;
      20'h0d470: out <= 12'h088;
      20'h0d471: out <= 12'h088;
      20'h0d472: out <= 12'h088;
      20'h0d473: out <= 12'h088;
      20'h0d474: out <= 12'h088;
      20'h0d475: out <= 12'h088;
      20'h0d476: out <= 12'h088;
      20'h0d477: out <= 12'h088;
      20'h0d478: out <= 12'h088;
      20'h0d479: out <= 12'h088;
      20'h0d47a: out <= 12'h088;
      20'h0d47b: out <= 12'h088;
      20'h0d47c: out <= 12'h088;
      20'h0d47d: out <= 12'h088;
      20'h0d47e: out <= 12'h088;
      20'h0d47f: out <= 12'h088;
      20'h0d480: out <= 12'h088;
      20'h0d481: out <= 12'h088;
      20'h0d482: out <= 12'h088;
      20'h0d483: out <= 12'h088;
      20'h0d484: out <= 12'h088;
      20'h0d485: out <= 12'h088;
      20'h0d486: out <= 12'h088;
      20'h0d487: out <= 12'h088;
      20'h0d488: out <= 12'h088;
      20'h0d489: out <= 12'h088;
      20'h0d48a: out <= 12'h088;
      20'h0d48b: out <= 12'h088;
      20'h0d48c: out <= 12'h088;
      20'h0d48d: out <= 12'h088;
      20'h0d48e: out <= 12'h088;
      20'h0d48f: out <= 12'h088;
      20'h0d490: out <= 12'h088;
      20'h0d491: out <= 12'h088;
      20'h0d492: out <= 12'h088;
      20'h0d493: out <= 12'h088;
      20'h0d494: out <= 12'h088;
      20'h0d495: out <= 12'h088;
      20'h0d496: out <= 12'h088;
      20'h0d497: out <= 12'h088;
      20'h0d498: out <= 12'h088;
      20'h0d499: out <= 12'hfff;
      20'h0d49a: out <= 12'hfff;
      20'h0d49b: out <= 12'hfff;
      20'h0d49c: out <= 12'hfff;
      20'h0d49d: out <= 12'h16d;
      20'h0d49e: out <= 12'h16d;
      20'h0d49f: out <= 12'h000;
      20'h0d4a0: out <= 12'h000;
      20'h0d4a1: out <= 12'h660;
      20'h0d4a2: out <= 12'h660;
      20'h0d4a3: out <= 12'hee9;
      20'h0d4a4: out <= 12'hee9;
      20'h0d4a5: out <= 12'hee9;
      20'h0d4a6: out <= 12'hee9;
      20'h0d4a7: out <= 12'hee9;
      20'h0d4a8: out <= 12'hee9;
      20'h0d4a9: out <= 12'hee9;
      20'h0d4aa: out <= 12'hee9;
      20'h0d4ab: out <= 12'hee9;
      20'h0d4ac: out <= 12'hee9;
      20'h0d4ad: out <= 12'h660;
      20'h0d4ae: out <= 12'h660;
      20'h0d4af: out <= 12'h000;
      20'h0d4b0: out <= 12'h603;
      20'h0d4b1: out <= 12'h603;
      20'h0d4b2: out <= 12'h603;
      20'h0d4b3: out <= 12'h603;
      20'h0d4b4: out <= 12'h603;
      20'h0d4b5: out <= 12'h603;
      20'h0d4b6: out <= 12'h603;
      20'h0d4b7: out <= 12'h603;
      20'h0d4b8: out <= 12'h603;
      20'h0d4b9: out <= 12'h603;
      20'h0d4ba: out <= 12'h603;
      20'h0d4bb: out <= 12'h603;
      20'h0d4bc: out <= 12'h603;
      20'h0d4bd: out <= 12'h603;
      20'h0d4be: out <= 12'h603;
      20'h0d4bf: out <= 12'h603;
      20'h0d4c0: out <= 12'h603;
      20'h0d4c1: out <= 12'h603;
      20'h0d4c2: out <= 12'h603;
      20'h0d4c3: out <= 12'h603;
      20'h0d4c4: out <= 12'h603;
      20'h0d4c5: out <= 12'h603;
      20'h0d4c6: out <= 12'h603;
      20'h0d4c7: out <= 12'h603;
      20'h0d4c8: out <= 12'h603;
      20'h0d4c9: out <= 12'h603;
      20'h0d4ca: out <= 12'h603;
      20'h0d4cb: out <= 12'h603;
      20'h0d4cc: out <= 12'h603;
      20'h0d4cd: out <= 12'h603;
      20'h0d4ce: out <= 12'h603;
      20'h0d4cf: out <= 12'h603;
      20'h0d4d0: out <= 12'h603;
      20'h0d4d1: out <= 12'h603;
      20'h0d4d2: out <= 12'h603;
      20'h0d4d3: out <= 12'h603;
      20'h0d4d4: out <= 12'h603;
      20'h0d4d5: out <= 12'h603;
      20'h0d4d6: out <= 12'h603;
      20'h0d4d7: out <= 12'h603;
      20'h0d4d8: out <= 12'h603;
      20'h0d4d9: out <= 12'h603;
      20'h0d4da: out <= 12'h603;
      20'h0d4db: out <= 12'h603;
      20'h0d4dc: out <= 12'h603;
      20'h0d4dd: out <= 12'h603;
      20'h0d4de: out <= 12'h603;
      20'h0d4df: out <= 12'h603;
      20'h0d4e0: out <= 12'h603;
      20'h0d4e1: out <= 12'h603;
      20'h0d4e2: out <= 12'h603;
      20'h0d4e3: out <= 12'h603;
      20'h0d4e4: out <= 12'h603;
      20'h0d4e5: out <= 12'h603;
      20'h0d4e6: out <= 12'h603;
      20'h0d4e7: out <= 12'h603;
      20'h0d4e8: out <= 12'h603;
      20'h0d4e9: out <= 12'h603;
      20'h0d4ea: out <= 12'h603;
      20'h0d4eb: out <= 12'h603;
      20'h0d4ec: out <= 12'h603;
      20'h0d4ed: out <= 12'h603;
      20'h0d4ee: out <= 12'h603;
      20'h0d4ef: out <= 12'h603;
      20'h0d4f0: out <= 12'h603;
      20'h0d4f1: out <= 12'h603;
      20'h0d4f2: out <= 12'h603;
      20'h0d4f3: out <= 12'h603;
      20'h0d4f4: out <= 12'h603;
      20'h0d4f5: out <= 12'h603;
      20'h0d4f6: out <= 12'h603;
      20'h0d4f7: out <= 12'h603;
      20'h0d4f8: out <= 12'h603;
      20'h0d4f9: out <= 12'h603;
      20'h0d4fa: out <= 12'h603;
      20'h0d4fb: out <= 12'h603;
      20'h0d4fc: out <= 12'h603;
      20'h0d4fd: out <= 12'h603;
      20'h0d4fe: out <= 12'h603;
      20'h0d4ff: out <= 12'h603;
      20'h0d500: out <= 12'h603;
      20'h0d501: out <= 12'h603;
      20'h0d502: out <= 12'h603;
      20'h0d503: out <= 12'h603;
      20'h0d504: out <= 12'h603;
      20'h0d505: out <= 12'h603;
      20'h0d506: out <= 12'h603;
      20'h0d507: out <= 12'h603;
      20'h0d508: out <= 12'hee9;
      20'h0d509: out <= 12'hf87;
      20'h0d50a: out <= 12'hee9;
      20'h0d50b: out <= 12'hee9;
      20'h0d50c: out <= 12'hee9;
      20'h0d50d: out <= 12'hb27;
      20'h0d50e: out <= 12'hf87;
      20'h0d50f: out <= 12'hb27;
      20'h0d510: out <= 12'h000;
      20'h0d511: out <= 12'h000;
      20'h0d512: out <= 12'h000;
      20'h0d513: out <= 12'h000;
      20'h0d514: out <= 12'h000;
      20'h0d515: out <= 12'h000;
      20'h0d516: out <= 12'h000;
      20'h0d517: out <= 12'h000;
      20'h0d518: out <= 12'hbbb;
      20'h0d519: out <= 12'hbbb;
      20'h0d51a: out <= 12'h000;
      20'h0d51b: out <= 12'h000;
      20'h0d51c: out <= 12'h000;
      20'h0d51d: out <= 12'h000;
      20'h0d51e: out <= 12'hbbb;
      20'h0d51f: out <= 12'hbbb;
      20'h0d520: out <= 12'h000;
      20'h0d521: out <= 12'h000;
      20'h0d522: out <= 12'hbbb;
      20'h0d523: out <= 12'hbbb;
      20'h0d524: out <= 12'h000;
      20'h0d525: out <= 12'hbbb;
      20'h0d526: out <= 12'hbbb;
      20'h0d527: out <= 12'h000;
      20'h0d528: out <= 12'h000;
      20'h0d529: out <= 12'h000;
      20'h0d52a: out <= 12'h000;
      20'h0d52b: out <= 12'hbbb;
      20'h0d52c: out <= 12'hbbb;
      20'h0d52d: out <= 12'h000;
      20'h0d52e: out <= 12'hbbb;
      20'h0d52f: out <= 12'hbbb;
      20'h0d530: out <= 12'h000;
      20'h0d531: out <= 12'hbbb;
      20'h0d532: out <= 12'hbbb;
      20'h0d533: out <= 12'h000;
      20'h0d534: out <= 12'hbbb;
      20'h0d535: out <= 12'hbbb;
      20'h0d536: out <= 12'h000;
      20'h0d537: out <= 12'h000;
      20'h0d538: out <= 12'h000;
      20'h0d539: out <= 12'hbbb;
      20'h0d53a: out <= 12'hbbb;
      20'h0d53b: out <= 12'h000;
      20'h0d53c: out <= 12'h000;
      20'h0d53d: out <= 12'h000;
      20'h0d53e: out <= 12'h000;
      20'h0d53f: out <= 12'h000;
      20'h0d540: out <= 12'h000;
      20'h0d541: out <= 12'h000;
      20'h0d542: out <= 12'h000;
      20'h0d543: out <= 12'h000;
      20'h0d544: out <= 12'h000;
      20'h0d545: out <= 12'h000;
      20'h0d546: out <= 12'h000;
      20'h0d547: out <= 12'h000;
      20'h0d548: out <= 12'h000;
      20'h0d549: out <= 12'h72f;
      20'h0d54a: out <= 12'hfff;
      20'h0d54b: out <= 12'hfff;
      20'h0d54c: out <= 12'hfff;
      20'h0d54d: out <= 12'hfff;
      20'h0d54e: out <= 12'h72f;
      20'h0d54f: out <= 12'h72f;
      20'h0d550: out <= 12'h72f;
      20'h0d551: out <= 12'h72f;
      20'h0d552: out <= 12'hfff;
      20'h0d553: out <= 12'hfff;
      20'h0d554: out <= 12'hfff;
      20'h0d555: out <= 12'hfff;
      20'h0d556: out <= 12'h72f;
      20'h0d557: out <= 12'h000;
      20'h0d558: out <= 12'h000;
      20'h0d559: out <= 12'h666;
      20'h0d55a: out <= 12'hfff;
      20'h0d55b: out <= 12'hfff;
      20'h0d55c: out <= 12'hfff;
      20'h0d55d: out <= 12'hfff;
      20'h0d55e: out <= 12'hfff;
      20'h0d55f: out <= 12'hfff;
      20'h0d560: out <= 12'h666;
      20'h0d561: out <= 12'h666;
      20'h0d562: out <= 12'h666;
      20'h0d563: out <= 12'hfff;
      20'h0d564: out <= 12'hfff;
      20'h0d565: out <= 12'hfff;
      20'h0d566: out <= 12'h666;
      20'h0d567: out <= 12'h000;
      20'h0d568: out <= 12'h000;
      20'h0d569: out <= 12'h660;
      20'h0d56a: out <= 12'hee9;
      20'h0d56b: out <= 12'hee9;
      20'h0d56c: out <= 12'hee9;
      20'h0d56d: out <= 12'hee9;
      20'h0d56e: out <= 12'h660;
      20'h0d56f: out <= 12'h660;
      20'h0d570: out <= 12'hbb0;
      20'h0d571: out <= 12'hbb0;
      20'h0d572: out <= 12'hee9;
      20'h0d573: out <= 12'hee9;
      20'h0d574: out <= 12'hee9;
      20'h0d575: out <= 12'hee9;
      20'h0d576: out <= 12'h660;
      20'h0d577: out <= 12'h000;
      20'h0d578: out <= 12'h000;
      20'h0d579: out <= 12'h16d;
      20'h0d57a: out <= 12'hfff;
      20'h0d57b: out <= 12'hfff;
      20'h0d57c: out <= 12'h6af;
      20'h0d57d: out <= 12'h16d;
      20'h0d57e: out <= 12'h16d;
      20'h0d57f: out <= 12'h16d;
      20'h0d580: out <= 12'h16d;
      20'h0d581: out <= 12'h16d;
      20'h0d582: out <= 12'h16d;
      20'h0d583: out <= 12'hfff;
      20'h0d584: out <= 12'hfff;
      20'h0d585: out <= 12'hfff;
      20'h0d586: out <= 12'h16d;
      20'h0d587: out <= 12'h000;
      20'h0d588: out <= 12'h000;
      20'h0d589: out <= 12'h72f;
      20'h0d58a: out <= 12'hfff;
      20'h0d58b: out <= 12'hfff;
      20'h0d58c: out <= 12'hfff;
      20'h0d58d: out <= 12'hfff;
      20'h0d58e: out <= 12'hfff;
      20'h0d58f: out <= 12'hfff;
      20'h0d590: out <= 12'hfff;
      20'h0d591: out <= 12'hfff;
      20'h0d592: out <= 12'hfff;
      20'h0d593: out <= 12'hfff;
      20'h0d594: out <= 12'hfff;
      20'h0d595: out <= 12'hfff;
      20'h0d596: out <= 12'h72f;
      20'h0d597: out <= 12'h000;
      20'h0d598: out <= 12'h000;
      20'h0d599: out <= 12'h666;
      20'h0d59a: out <= 12'hfff;
      20'h0d59b: out <= 12'hfff;
      20'h0d59c: out <= 12'hfff;
      20'h0d59d: out <= 12'h666;
      20'h0d59e: out <= 12'hbbb;
      20'h0d59f: out <= 12'hfff;
      20'h0d5a0: out <= 12'hfff;
      20'h0d5a1: out <= 12'hfff;
      20'h0d5a2: out <= 12'hfff;
      20'h0d5a3: out <= 12'hfff;
      20'h0d5a4: out <= 12'hfff;
      20'h0d5a5: out <= 12'hfff;
      20'h0d5a6: out <= 12'h666;
      20'h0d5a7: out <= 12'h000;
      20'h0d5a8: out <= 12'h000;
      20'h0d5a9: out <= 12'h16d;
      20'h0d5aa: out <= 12'hfff;
      20'h0d5ab: out <= 12'hfff;
      20'h0d5ac: out <= 12'hfff;
      20'h0d5ad: out <= 12'hfff;
      20'h0d5ae: out <= 12'hfff;
      20'h0d5af: out <= 12'h6af;
      20'h0d5b0: out <= 12'h16d;
      20'h0d5b1: out <= 12'hfff;
      20'h0d5b2: out <= 12'hfff;
      20'h0d5b3: out <= 12'hfff;
      20'h0d5b4: out <= 12'hfff;
      20'h0d5b5: out <= 12'hfff;
      20'h0d5b6: out <= 12'h16d;
      20'h0d5b7: out <= 12'h000;
      20'h0d5b8: out <= 12'h000;
      20'h0d5b9: out <= 12'h660;
      20'h0d5ba: out <= 12'hee9;
      20'h0d5bb: out <= 12'hee9;
      20'h0d5bc: out <= 12'hee9;
      20'h0d5bd: out <= 12'hee9;
      20'h0d5be: out <= 12'h660;
      20'h0d5bf: out <= 12'h660;
      20'h0d5c0: out <= 12'h660;
      20'h0d5c1: out <= 12'h660;
      20'h0d5c2: out <= 12'hee9;
      20'h0d5c3: out <= 12'hee9;
      20'h0d5c4: out <= 12'hee9;
      20'h0d5c5: out <= 12'hee9;
      20'h0d5c6: out <= 12'h660;
      20'h0d5c7: out <= 12'h000;
      20'h0d5c8: out <= 12'h603;
      20'h0d5c9: out <= 12'h603;
      20'h0d5ca: out <= 12'h603;
      20'h0d5cb: out <= 12'h603;
      20'h0d5cc: out <= 12'h603;
      20'h0d5cd: out <= 12'h603;
      20'h0d5ce: out <= 12'h603;
      20'h0d5cf: out <= 12'h603;
      20'h0d5d0: out <= 12'h603;
      20'h0d5d1: out <= 12'h603;
      20'h0d5d2: out <= 12'h603;
      20'h0d5d3: out <= 12'h603;
      20'h0d5d4: out <= 12'h603;
      20'h0d5d5: out <= 12'h603;
      20'h0d5d6: out <= 12'h603;
      20'h0d5d7: out <= 12'h603;
      20'h0d5d8: out <= 12'h603;
      20'h0d5d9: out <= 12'h603;
      20'h0d5da: out <= 12'h603;
      20'h0d5db: out <= 12'h603;
      20'h0d5dc: out <= 12'h603;
      20'h0d5dd: out <= 12'h603;
      20'h0d5de: out <= 12'h603;
      20'h0d5df: out <= 12'h603;
      20'h0d5e0: out <= 12'h603;
      20'h0d5e1: out <= 12'h603;
      20'h0d5e2: out <= 12'h603;
      20'h0d5e3: out <= 12'h603;
      20'h0d5e4: out <= 12'h603;
      20'h0d5e5: out <= 12'h603;
      20'h0d5e6: out <= 12'h603;
      20'h0d5e7: out <= 12'h603;
      20'h0d5e8: out <= 12'h603;
      20'h0d5e9: out <= 12'h603;
      20'h0d5ea: out <= 12'h603;
      20'h0d5eb: out <= 12'h603;
      20'h0d5ec: out <= 12'h603;
      20'h0d5ed: out <= 12'h603;
      20'h0d5ee: out <= 12'h603;
      20'h0d5ef: out <= 12'h603;
      20'h0d5f0: out <= 12'h603;
      20'h0d5f1: out <= 12'h603;
      20'h0d5f2: out <= 12'h603;
      20'h0d5f3: out <= 12'h603;
      20'h0d5f4: out <= 12'h603;
      20'h0d5f5: out <= 12'h603;
      20'h0d5f6: out <= 12'h603;
      20'h0d5f7: out <= 12'h603;
      20'h0d5f8: out <= 12'h603;
      20'h0d5f9: out <= 12'h603;
      20'h0d5fa: out <= 12'h603;
      20'h0d5fb: out <= 12'h603;
      20'h0d5fc: out <= 12'h603;
      20'h0d5fd: out <= 12'h603;
      20'h0d5fe: out <= 12'h603;
      20'h0d5ff: out <= 12'h603;
      20'h0d600: out <= 12'h603;
      20'h0d601: out <= 12'h603;
      20'h0d602: out <= 12'h603;
      20'h0d603: out <= 12'h603;
      20'h0d604: out <= 12'h603;
      20'h0d605: out <= 12'h603;
      20'h0d606: out <= 12'h603;
      20'h0d607: out <= 12'h603;
      20'h0d608: out <= 12'h603;
      20'h0d609: out <= 12'h603;
      20'h0d60a: out <= 12'h603;
      20'h0d60b: out <= 12'h603;
      20'h0d60c: out <= 12'h603;
      20'h0d60d: out <= 12'h603;
      20'h0d60e: out <= 12'h603;
      20'h0d60f: out <= 12'h603;
      20'h0d610: out <= 12'h603;
      20'h0d611: out <= 12'h603;
      20'h0d612: out <= 12'h603;
      20'h0d613: out <= 12'h603;
      20'h0d614: out <= 12'h603;
      20'h0d615: out <= 12'h603;
      20'h0d616: out <= 12'h603;
      20'h0d617: out <= 12'h603;
      20'h0d618: out <= 12'h603;
      20'h0d619: out <= 12'h603;
      20'h0d61a: out <= 12'h603;
      20'h0d61b: out <= 12'h603;
      20'h0d61c: out <= 12'h603;
      20'h0d61d: out <= 12'h603;
      20'h0d61e: out <= 12'h603;
      20'h0d61f: out <= 12'h603;
      20'h0d620: out <= 12'hee9;
      20'h0d621: out <= 12'hf87;
      20'h0d622: out <= 12'hee9;
      20'h0d623: out <= 12'hf87;
      20'h0d624: out <= 12'hf87;
      20'h0d625: out <= 12'hb27;
      20'h0d626: out <= 12'hf87;
      20'h0d627: out <= 12'hb27;
      20'h0d628: out <= 12'h000;
      20'h0d629: out <= 12'h000;
      20'h0d62a: out <= 12'h000;
      20'h0d62b: out <= 12'h000;
      20'h0d62c: out <= 12'h000;
      20'h0d62d: out <= 12'h000;
      20'h0d62e: out <= 12'h000;
      20'h0d62f: out <= 12'h000;
      20'h0d630: out <= 12'hbbb;
      20'h0d631: out <= 12'hbbb;
      20'h0d632: out <= 12'hbbb;
      20'h0d633: out <= 12'hbbb;
      20'h0d634: out <= 12'h000;
      20'h0d635: out <= 12'h000;
      20'h0d636: out <= 12'hbbb;
      20'h0d637: out <= 12'hbbb;
      20'h0d638: out <= 12'h000;
      20'h0d639: out <= 12'h000;
      20'h0d63a: out <= 12'hbbb;
      20'h0d63b: out <= 12'hbbb;
      20'h0d63c: out <= 12'h000;
      20'h0d63d: out <= 12'hbbb;
      20'h0d63e: out <= 12'hbbb;
      20'h0d63f: out <= 12'hbbb;
      20'h0d640: out <= 12'hbbb;
      20'h0d641: out <= 12'h000;
      20'h0d642: out <= 12'h000;
      20'h0d643: out <= 12'hbbb;
      20'h0d644: out <= 12'hbbb;
      20'h0d645: out <= 12'h000;
      20'h0d646: out <= 12'hbbb;
      20'h0d647: out <= 12'hbbb;
      20'h0d648: out <= 12'h000;
      20'h0d649: out <= 12'hbbb;
      20'h0d64a: out <= 12'hbbb;
      20'h0d64b: out <= 12'h000;
      20'h0d64c: out <= 12'h000;
      20'h0d64d: out <= 12'hbbb;
      20'h0d64e: out <= 12'hbbb;
      20'h0d64f: out <= 12'hbbb;
      20'h0d650: out <= 12'hbbb;
      20'h0d651: out <= 12'hbbb;
      20'h0d652: out <= 12'h000;
      20'h0d653: out <= 12'h000;
      20'h0d654: out <= 12'h000;
      20'h0d655: out <= 12'h000;
      20'h0d656: out <= 12'h000;
      20'h0d657: out <= 12'h000;
      20'h0d658: out <= 12'h000;
      20'h0d659: out <= 12'h000;
      20'h0d65a: out <= 12'h000;
      20'h0d65b: out <= 12'h000;
      20'h0d65c: out <= 12'h000;
      20'h0d65d: out <= 12'h000;
      20'h0d65e: out <= 12'h000;
      20'h0d65f: out <= 12'h000;
      20'h0d660: out <= 12'h000;
      20'h0d661: out <= 12'h72f;
      20'h0d662: out <= 12'hfff;
      20'h0d663: out <= 12'hfff;
      20'h0d664: out <= 12'hc7f;
      20'h0d665: out <= 12'h72f;
      20'h0d666: out <= 12'hc7f;
      20'h0d667: out <= 12'hc7f;
      20'h0d668: out <= 12'hc7f;
      20'h0d669: out <= 12'hc7f;
      20'h0d66a: out <= 12'h72f;
      20'h0d66b: out <= 12'hc7f;
      20'h0d66c: out <= 12'hfff;
      20'h0d66d: out <= 12'hfff;
      20'h0d66e: out <= 12'h72f;
      20'h0d66f: out <= 12'h000;
      20'h0d670: out <= 12'h000;
      20'h0d671: out <= 12'h666;
      20'h0d672: out <= 12'hfff;
      20'h0d673: out <= 12'hfff;
      20'h0d674: out <= 12'hfff;
      20'h0d675: out <= 12'hfff;
      20'h0d676: out <= 12'hfff;
      20'h0d677: out <= 12'h666;
      20'h0d678: out <= 12'hfff;
      20'h0d679: out <= 12'hfff;
      20'h0d67a: out <= 12'hfff;
      20'h0d67b: out <= 12'hfff;
      20'h0d67c: out <= 12'hfff;
      20'h0d67d: out <= 12'hfff;
      20'h0d67e: out <= 12'h666;
      20'h0d67f: out <= 12'h000;
      20'h0d680: out <= 12'h000;
      20'h0d681: out <= 12'h660;
      20'h0d682: out <= 12'hee9;
      20'h0d683: out <= 12'hbb0;
      20'h0d684: out <= 12'hbb0;
      20'h0d685: out <= 12'hee9;
      20'h0d686: out <= 12'hee9;
      20'h0d687: out <= 12'h660;
      20'h0d688: out <= 12'hbb0;
      20'h0d689: out <= 12'hee9;
      20'h0d68a: out <= 12'hee9;
      20'h0d68b: out <= 12'hbb0;
      20'h0d68c: out <= 12'hbb0;
      20'h0d68d: out <= 12'hee9;
      20'h0d68e: out <= 12'h660;
      20'h0d68f: out <= 12'h000;
      20'h0d690: out <= 12'h000;
      20'h0d691: out <= 12'h16d;
      20'h0d692: out <= 12'hfff;
      20'h0d693: out <= 12'hfff;
      20'h0d694: out <= 12'h6af;
      20'h0d695: out <= 12'h16d;
      20'h0d696: out <= 12'h16d;
      20'h0d697: out <= 12'hfff;
      20'h0d698: out <= 12'hfff;
      20'h0d699: out <= 12'h6af;
      20'h0d69a: out <= 12'h16d;
      20'h0d69b: out <= 12'h16d;
      20'h0d69c: out <= 12'hfff;
      20'h0d69d: out <= 12'hfff;
      20'h0d69e: out <= 12'h16d;
      20'h0d69f: out <= 12'h000;
      20'h0d6a0: out <= 12'h000;
      20'h0d6a1: out <= 12'h72f;
      20'h0d6a2: out <= 12'hfff;
      20'h0d6a3: out <= 12'h72f;
      20'h0d6a4: out <= 12'hfff;
      20'h0d6a5: out <= 12'hfff;
      20'h0d6a6: out <= 12'hfff;
      20'h0d6a7: out <= 12'hfff;
      20'h0d6a8: out <= 12'hfff;
      20'h0d6a9: out <= 12'hfff;
      20'h0d6aa: out <= 12'hfff;
      20'h0d6ab: out <= 12'hfff;
      20'h0d6ac: out <= 12'h72f;
      20'h0d6ad: out <= 12'hfff;
      20'h0d6ae: out <= 12'h72f;
      20'h0d6af: out <= 12'h000;
      20'h0d6b0: out <= 12'h000;
      20'h0d6b1: out <= 12'h666;
      20'h0d6b2: out <= 12'hfff;
      20'h0d6b3: out <= 12'hfff;
      20'h0d6b4: out <= 12'hfff;
      20'h0d6b5: out <= 12'h666;
      20'h0d6b6: out <= 12'hbbb;
      20'h0d6b7: out <= 12'h666;
      20'h0d6b8: out <= 12'hfff;
      20'h0d6b9: out <= 12'hfff;
      20'h0d6ba: out <= 12'hfff;
      20'h0d6bb: out <= 12'hfff;
      20'h0d6bc: out <= 12'hfff;
      20'h0d6bd: out <= 12'hfff;
      20'h0d6be: out <= 12'h666;
      20'h0d6bf: out <= 12'h000;
      20'h0d6c0: out <= 12'h000;
      20'h0d6c1: out <= 12'h16d;
      20'h0d6c2: out <= 12'hfff;
      20'h0d6c3: out <= 12'hfff;
      20'h0d6c4: out <= 12'hfff;
      20'h0d6c5: out <= 12'hfff;
      20'h0d6c6: out <= 12'h6af;
      20'h0d6c7: out <= 12'h16d;
      20'h0d6c8: out <= 12'h6af;
      20'h0d6c9: out <= 12'h16d;
      20'h0d6ca: out <= 12'hfff;
      20'h0d6cb: out <= 12'hfff;
      20'h0d6cc: out <= 12'hfff;
      20'h0d6cd: out <= 12'hfff;
      20'h0d6ce: out <= 12'h16d;
      20'h0d6cf: out <= 12'h000;
      20'h0d6d0: out <= 12'h000;
      20'h0d6d1: out <= 12'h660;
      20'h0d6d2: out <= 12'hee9;
      20'h0d6d3: out <= 12'hee9;
      20'h0d6d4: out <= 12'hee9;
      20'h0d6d5: out <= 12'h660;
      20'h0d6d6: out <= 12'hbb0;
      20'h0d6d7: out <= 12'hbb0;
      20'h0d6d8: out <= 12'hbb0;
      20'h0d6d9: out <= 12'hbb0;
      20'h0d6da: out <= 12'h660;
      20'h0d6db: out <= 12'hee9;
      20'h0d6dc: out <= 12'hee9;
      20'h0d6dd: out <= 12'hee9;
      20'h0d6de: out <= 12'h660;
      20'h0d6df: out <= 12'h000;
      20'h0d6e0: out <= 12'h603;
      20'h0d6e1: out <= 12'h603;
      20'h0d6e2: out <= 12'h603;
      20'h0d6e3: out <= 12'h603;
      20'h0d6e4: out <= 12'h603;
      20'h0d6e5: out <= 12'h603;
      20'h0d6e6: out <= 12'h603;
      20'h0d6e7: out <= 12'h603;
      20'h0d6e8: out <= 12'h603;
      20'h0d6e9: out <= 12'h603;
      20'h0d6ea: out <= 12'h603;
      20'h0d6eb: out <= 12'h603;
      20'h0d6ec: out <= 12'h603;
      20'h0d6ed: out <= 12'h603;
      20'h0d6ee: out <= 12'h603;
      20'h0d6ef: out <= 12'h603;
      20'h0d6f0: out <= 12'h603;
      20'h0d6f1: out <= 12'h603;
      20'h0d6f2: out <= 12'h603;
      20'h0d6f3: out <= 12'h603;
      20'h0d6f4: out <= 12'h603;
      20'h0d6f5: out <= 12'h603;
      20'h0d6f6: out <= 12'h603;
      20'h0d6f7: out <= 12'h603;
      20'h0d6f8: out <= 12'h603;
      20'h0d6f9: out <= 12'h603;
      20'h0d6fa: out <= 12'h603;
      20'h0d6fb: out <= 12'h603;
      20'h0d6fc: out <= 12'h603;
      20'h0d6fd: out <= 12'h603;
      20'h0d6fe: out <= 12'h603;
      20'h0d6ff: out <= 12'h603;
      20'h0d700: out <= 12'h603;
      20'h0d701: out <= 12'h603;
      20'h0d702: out <= 12'h603;
      20'h0d703: out <= 12'h603;
      20'h0d704: out <= 12'h603;
      20'h0d705: out <= 12'h603;
      20'h0d706: out <= 12'h603;
      20'h0d707: out <= 12'h603;
      20'h0d708: out <= 12'h603;
      20'h0d709: out <= 12'h603;
      20'h0d70a: out <= 12'h603;
      20'h0d70b: out <= 12'h603;
      20'h0d70c: out <= 12'h603;
      20'h0d70d: out <= 12'h603;
      20'h0d70e: out <= 12'h603;
      20'h0d70f: out <= 12'h603;
      20'h0d710: out <= 12'h603;
      20'h0d711: out <= 12'h603;
      20'h0d712: out <= 12'h603;
      20'h0d713: out <= 12'h603;
      20'h0d714: out <= 12'h603;
      20'h0d715: out <= 12'h603;
      20'h0d716: out <= 12'h603;
      20'h0d717: out <= 12'h603;
      20'h0d718: out <= 12'h603;
      20'h0d719: out <= 12'h603;
      20'h0d71a: out <= 12'h603;
      20'h0d71b: out <= 12'h603;
      20'h0d71c: out <= 12'h603;
      20'h0d71d: out <= 12'h603;
      20'h0d71e: out <= 12'h603;
      20'h0d71f: out <= 12'h603;
      20'h0d720: out <= 12'h603;
      20'h0d721: out <= 12'h603;
      20'h0d722: out <= 12'h603;
      20'h0d723: out <= 12'h603;
      20'h0d724: out <= 12'h603;
      20'h0d725: out <= 12'h603;
      20'h0d726: out <= 12'h603;
      20'h0d727: out <= 12'h603;
      20'h0d728: out <= 12'h603;
      20'h0d729: out <= 12'h603;
      20'h0d72a: out <= 12'h603;
      20'h0d72b: out <= 12'h603;
      20'h0d72c: out <= 12'h603;
      20'h0d72d: out <= 12'h603;
      20'h0d72e: out <= 12'h603;
      20'h0d72f: out <= 12'h603;
      20'h0d730: out <= 12'h603;
      20'h0d731: out <= 12'h603;
      20'h0d732: out <= 12'h603;
      20'h0d733: out <= 12'h603;
      20'h0d734: out <= 12'h603;
      20'h0d735: out <= 12'h603;
      20'h0d736: out <= 12'h603;
      20'h0d737: out <= 12'h603;
      20'h0d738: out <= 12'hee9;
      20'h0d739: out <= 12'hf87;
      20'h0d73a: out <= 12'hee9;
      20'h0d73b: out <= 12'hf87;
      20'h0d73c: out <= 12'hf87;
      20'h0d73d: out <= 12'hb27;
      20'h0d73e: out <= 12'hf87;
      20'h0d73f: out <= 12'hb27;
      20'h0d740: out <= 12'h000;
      20'h0d741: out <= 12'h000;
      20'h0d742: out <= 12'h000;
      20'h0d743: out <= 12'h000;
      20'h0d744: out <= 12'h000;
      20'h0d745: out <= 12'h000;
      20'h0d746: out <= 12'h000;
      20'h0d747: out <= 12'h000;
      20'h0d748: out <= 12'hbbb;
      20'h0d749: out <= 12'hbbb;
      20'h0d74a: out <= 12'h000;
      20'h0d74b: out <= 12'h000;
      20'h0d74c: out <= 12'h000;
      20'h0d74d: out <= 12'h000;
      20'h0d74e: out <= 12'hbbb;
      20'h0d74f: out <= 12'hbbb;
      20'h0d750: out <= 12'h000;
      20'h0d751: out <= 12'h000;
      20'h0d752: out <= 12'hbbb;
      20'h0d753: out <= 12'hbbb;
      20'h0d754: out <= 12'h000;
      20'h0d755: out <= 12'hbbb;
      20'h0d756: out <= 12'hbbb;
      20'h0d757: out <= 12'h000;
      20'h0d758: out <= 12'h000;
      20'h0d759: out <= 12'h000;
      20'h0d75a: out <= 12'h000;
      20'h0d75b: out <= 12'hbbb;
      20'h0d75c: out <= 12'hbbb;
      20'h0d75d: out <= 12'h000;
      20'h0d75e: out <= 12'hbbb;
      20'h0d75f: out <= 12'hbbb;
      20'h0d760: out <= 12'h000;
      20'h0d761: out <= 12'hbbb;
      20'h0d762: out <= 12'hbbb;
      20'h0d763: out <= 12'h000;
      20'h0d764: out <= 12'h000;
      20'h0d765: out <= 12'h000;
      20'h0d766: out <= 12'hbbb;
      20'h0d767: out <= 12'hbbb;
      20'h0d768: out <= 12'hbbb;
      20'h0d769: out <= 12'h000;
      20'h0d76a: out <= 12'h000;
      20'h0d76b: out <= 12'h000;
      20'h0d76c: out <= 12'h000;
      20'h0d76d: out <= 12'h000;
      20'h0d76e: out <= 12'h000;
      20'h0d76f: out <= 12'h000;
      20'h0d770: out <= 12'h000;
      20'h0d771: out <= 12'h000;
      20'h0d772: out <= 12'h000;
      20'h0d773: out <= 12'h000;
      20'h0d774: out <= 12'h000;
      20'h0d775: out <= 12'h000;
      20'h0d776: out <= 12'h000;
      20'h0d777: out <= 12'h000;
      20'h0d778: out <= 12'h000;
      20'h0d779: out <= 12'hc7f;
      20'h0d77a: out <= 12'hfff;
      20'h0d77b: out <= 12'hfff;
      20'h0d77c: out <= 12'h72f;
      20'h0d77d: out <= 12'hc7f;
      20'h0d77e: out <= 12'hfff;
      20'h0d77f: out <= 12'hfff;
      20'h0d780: out <= 12'h72f;
      20'h0d781: out <= 12'hfff;
      20'h0d782: out <= 12'hc7f;
      20'h0d783: out <= 12'h72f;
      20'h0d784: out <= 12'hfff;
      20'h0d785: out <= 12'hfff;
      20'h0d786: out <= 12'hc7f;
      20'h0d787: out <= 12'h000;
      20'h0d788: out <= 12'h000;
      20'h0d789: out <= 12'hbbb;
      20'h0d78a: out <= 12'hfff;
      20'h0d78b: out <= 12'hfff;
      20'h0d78c: out <= 12'hfff;
      20'h0d78d: out <= 12'h666;
      20'h0d78e: out <= 12'h666;
      20'h0d78f: out <= 12'h666;
      20'h0d790: out <= 12'h666;
      20'h0d791: out <= 12'h666;
      20'h0d792: out <= 12'h666;
      20'h0d793: out <= 12'hfff;
      20'h0d794: out <= 12'hfff;
      20'h0d795: out <= 12'hfff;
      20'h0d796: out <= 12'hbbb;
      20'h0d797: out <= 12'h000;
      20'h0d798: out <= 12'h000;
      20'h0d799: out <= 12'hbb0;
      20'h0d79a: out <= 12'hee9;
      20'h0d79b: out <= 12'h660;
      20'h0d79c: out <= 12'h660;
      20'h0d79d: out <= 12'hee9;
      20'h0d79e: out <= 12'hee9;
      20'h0d79f: out <= 12'h660;
      20'h0d7a0: out <= 12'hbb0;
      20'h0d7a1: out <= 12'hee9;
      20'h0d7a2: out <= 12'hee9;
      20'h0d7a3: out <= 12'h660;
      20'h0d7a4: out <= 12'h660;
      20'h0d7a5: out <= 12'hee9;
      20'h0d7a6: out <= 12'hbb0;
      20'h0d7a7: out <= 12'h000;
      20'h0d7a8: out <= 12'h000;
      20'h0d7a9: out <= 12'h6af;
      20'h0d7aa: out <= 12'hfff;
      20'h0d7ab: out <= 12'hfff;
      20'h0d7ac: out <= 12'h6af;
      20'h0d7ad: out <= 12'h16d;
      20'h0d7ae: out <= 12'h16d;
      20'h0d7af: out <= 12'hfff;
      20'h0d7b0: out <= 12'hfff;
      20'h0d7b1: out <= 12'h6af;
      20'h0d7b2: out <= 12'h16d;
      20'h0d7b3: out <= 12'h16d;
      20'h0d7b4: out <= 12'hfff;
      20'h0d7b5: out <= 12'hfff;
      20'h0d7b6: out <= 12'h6af;
      20'h0d7b7: out <= 12'h000;
      20'h0d7b8: out <= 12'h000;
      20'h0d7b9: out <= 12'hc7f;
      20'h0d7ba: out <= 12'hfff;
      20'h0d7bb: out <= 12'h72f;
      20'h0d7bc: out <= 12'h72f;
      20'h0d7bd: out <= 12'hc7f;
      20'h0d7be: out <= 12'hc7f;
      20'h0d7bf: out <= 12'hc7f;
      20'h0d7c0: out <= 12'hc7f;
      20'h0d7c1: out <= 12'hc7f;
      20'h0d7c2: out <= 12'hc7f;
      20'h0d7c3: out <= 12'h72f;
      20'h0d7c4: out <= 12'h72f;
      20'h0d7c5: out <= 12'hfff;
      20'h0d7c6: out <= 12'hc7f;
      20'h0d7c7: out <= 12'h000;
      20'h0d7c8: out <= 12'h000;
      20'h0d7c9: out <= 12'hbbb;
      20'h0d7ca: out <= 12'hfff;
      20'h0d7cb: out <= 12'hfff;
      20'h0d7cc: out <= 12'hfff;
      20'h0d7cd: out <= 12'h666;
      20'h0d7ce: out <= 12'hbbb;
      20'h0d7cf: out <= 12'h666;
      20'h0d7d0: out <= 12'hbbb;
      20'h0d7d1: out <= 12'hfff;
      20'h0d7d2: out <= 12'hfff;
      20'h0d7d3: out <= 12'hfff;
      20'h0d7d4: out <= 12'hfff;
      20'h0d7d5: out <= 12'hfff;
      20'h0d7d6: out <= 12'hbbb;
      20'h0d7d7: out <= 12'h000;
      20'h0d7d8: out <= 12'h000;
      20'h0d7d9: out <= 12'h6af;
      20'h0d7da: out <= 12'hfff;
      20'h0d7db: out <= 12'hfff;
      20'h0d7dc: out <= 12'hfff;
      20'h0d7dd: out <= 12'h6af;
      20'h0d7de: out <= 12'h6af;
      20'h0d7df: out <= 12'h16d;
      20'h0d7e0: out <= 12'h6af;
      20'h0d7e1: out <= 12'h16d;
      20'h0d7e2: out <= 12'h16d;
      20'h0d7e3: out <= 12'hfff;
      20'h0d7e4: out <= 12'hfff;
      20'h0d7e5: out <= 12'hfff;
      20'h0d7e6: out <= 12'h6af;
      20'h0d7e7: out <= 12'h000;
      20'h0d7e8: out <= 12'h000;
      20'h0d7e9: out <= 12'hbb0;
      20'h0d7ea: out <= 12'hee9;
      20'h0d7eb: out <= 12'hee9;
      20'h0d7ec: out <= 12'h660;
      20'h0d7ed: out <= 12'hbb0;
      20'h0d7ee: out <= 12'hbb0;
      20'h0d7ef: out <= 12'hee9;
      20'h0d7f0: out <= 12'hee9;
      20'h0d7f1: out <= 12'hbb0;
      20'h0d7f2: out <= 12'hbb0;
      20'h0d7f3: out <= 12'h660;
      20'h0d7f4: out <= 12'hee9;
      20'h0d7f5: out <= 12'hee9;
      20'h0d7f6: out <= 12'hbb0;
      20'h0d7f7: out <= 12'h000;
      20'h0d7f8: out <= 12'h603;
      20'h0d7f9: out <= 12'h603;
      20'h0d7fa: out <= 12'h603;
      20'h0d7fb: out <= 12'h603;
      20'h0d7fc: out <= 12'h603;
      20'h0d7fd: out <= 12'h603;
      20'h0d7fe: out <= 12'h603;
      20'h0d7ff: out <= 12'h603;
      20'h0d800: out <= 12'h603;
      20'h0d801: out <= 12'h603;
      20'h0d802: out <= 12'h603;
      20'h0d803: out <= 12'h603;
      20'h0d804: out <= 12'h603;
      20'h0d805: out <= 12'h603;
      20'h0d806: out <= 12'h603;
      20'h0d807: out <= 12'h603;
      20'h0d808: out <= 12'h603;
      20'h0d809: out <= 12'h603;
      20'h0d80a: out <= 12'h603;
      20'h0d80b: out <= 12'h603;
      20'h0d80c: out <= 12'h603;
      20'h0d80d: out <= 12'h603;
      20'h0d80e: out <= 12'h603;
      20'h0d80f: out <= 12'h603;
      20'h0d810: out <= 12'h603;
      20'h0d811: out <= 12'h603;
      20'h0d812: out <= 12'h603;
      20'h0d813: out <= 12'h603;
      20'h0d814: out <= 12'h603;
      20'h0d815: out <= 12'h603;
      20'h0d816: out <= 12'h603;
      20'h0d817: out <= 12'h603;
      20'h0d818: out <= 12'h603;
      20'h0d819: out <= 12'h603;
      20'h0d81a: out <= 12'h603;
      20'h0d81b: out <= 12'h603;
      20'h0d81c: out <= 12'h603;
      20'h0d81d: out <= 12'h603;
      20'h0d81e: out <= 12'h603;
      20'h0d81f: out <= 12'h603;
      20'h0d820: out <= 12'h603;
      20'h0d821: out <= 12'h603;
      20'h0d822: out <= 12'h603;
      20'h0d823: out <= 12'h603;
      20'h0d824: out <= 12'h603;
      20'h0d825: out <= 12'h603;
      20'h0d826: out <= 12'h603;
      20'h0d827: out <= 12'h603;
      20'h0d828: out <= 12'h603;
      20'h0d829: out <= 12'h603;
      20'h0d82a: out <= 12'h603;
      20'h0d82b: out <= 12'h603;
      20'h0d82c: out <= 12'h603;
      20'h0d82d: out <= 12'h603;
      20'h0d82e: out <= 12'h603;
      20'h0d82f: out <= 12'h603;
      20'h0d830: out <= 12'h603;
      20'h0d831: out <= 12'h603;
      20'h0d832: out <= 12'h603;
      20'h0d833: out <= 12'h603;
      20'h0d834: out <= 12'h603;
      20'h0d835: out <= 12'h603;
      20'h0d836: out <= 12'h603;
      20'h0d837: out <= 12'h603;
      20'h0d838: out <= 12'h603;
      20'h0d839: out <= 12'h603;
      20'h0d83a: out <= 12'h603;
      20'h0d83b: out <= 12'h603;
      20'h0d83c: out <= 12'h603;
      20'h0d83d: out <= 12'h603;
      20'h0d83e: out <= 12'h603;
      20'h0d83f: out <= 12'h603;
      20'h0d840: out <= 12'h603;
      20'h0d841: out <= 12'h603;
      20'h0d842: out <= 12'h603;
      20'h0d843: out <= 12'h603;
      20'h0d844: out <= 12'h603;
      20'h0d845: out <= 12'h603;
      20'h0d846: out <= 12'h603;
      20'h0d847: out <= 12'h603;
      20'h0d848: out <= 12'h603;
      20'h0d849: out <= 12'h603;
      20'h0d84a: out <= 12'h603;
      20'h0d84b: out <= 12'h603;
      20'h0d84c: out <= 12'h603;
      20'h0d84d: out <= 12'h603;
      20'h0d84e: out <= 12'h603;
      20'h0d84f: out <= 12'h603;
      20'h0d850: out <= 12'hee9;
      20'h0d851: out <= 12'hf87;
      20'h0d852: out <= 12'hee9;
      20'h0d853: out <= 12'hb27;
      20'h0d854: out <= 12'hb27;
      20'h0d855: out <= 12'hb27;
      20'h0d856: out <= 12'hf87;
      20'h0d857: out <= 12'hb27;
      20'h0d858: out <= 12'h000;
      20'h0d859: out <= 12'h000;
      20'h0d85a: out <= 12'h000;
      20'h0d85b: out <= 12'h000;
      20'h0d85c: out <= 12'h000;
      20'h0d85d: out <= 12'h000;
      20'h0d85e: out <= 12'h000;
      20'h0d85f: out <= 12'h000;
      20'h0d860: out <= 12'hbbb;
      20'h0d861: out <= 12'hbbb;
      20'h0d862: out <= 12'h000;
      20'h0d863: out <= 12'h000;
      20'h0d864: out <= 12'h000;
      20'h0d865: out <= 12'h000;
      20'h0d866: out <= 12'hbbb;
      20'h0d867: out <= 12'hbbb;
      20'h0d868: out <= 12'h000;
      20'h0d869: out <= 12'h000;
      20'h0d86a: out <= 12'hbbb;
      20'h0d86b: out <= 12'hbbb;
      20'h0d86c: out <= 12'h000;
      20'h0d86d: out <= 12'hbbb;
      20'h0d86e: out <= 12'hbbb;
      20'h0d86f: out <= 12'h000;
      20'h0d870: out <= 12'h000;
      20'h0d871: out <= 12'h000;
      20'h0d872: out <= 12'h000;
      20'h0d873: out <= 12'hbbb;
      20'h0d874: out <= 12'hbbb;
      20'h0d875: out <= 12'h000;
      20'h0d876: out <= 12'hbbb;
      20'h0d877: out <= 12'hbbb;
      20'h0d878: out <= 12'h000;
      20'h0d879: out <= 12'hbbb;
      20'h0d87a: out <= 12'hbbb;
      20'h0d87b: out <= 12'h000;
      20'h0d87c: out <= 12'h000;
      20'h0d87d: out <= 12'h000;
      20'h0d87e: out <= 12'hbbb;
      20'h0d87f: out <= 12'hbbb;
      20'h0d880: out <= 12'hbbb;
      20'h0d881: out <= 12'h000;
      20'h0d882: out <= 12'h000;
      20'h0d883: out <= 12'h000;
      20'h0d884: out <= 12'h000;
      20'h0d885: out <= 12'h000;
      20'h0d886: out <= 12'h000;
      20'h0d887: out <= 12'h000;
      20'h0d888: out <= 12'h000;
      20'h0d889: out <= 12'h000;
      20'h0d88a: out <= 12'h000;
      20'h0d88b: out <= 12'h000;
      20'h0d88c: out <= 12'h000;
      20'h0d88d: out <= 12'h000;
      20'h0d88e: out <= 12'h000;
      20'h0d88f: out <= 12'h000;
      20'h0d890: out <= 12'h000;
      20'h0d891: out <= 12'hc7f;
      20'h0d892: out <= 12'hfff;
      20'h0d893: out <= 12'h72f;
      20'h0d894: out <= 12'hc7f;
      20'h0d895: out <= 12'hfff;
      20'h0d896: out <= 12'hfff;
      20'h0d897: out <= 12'hfff;
      20'h0d898: out <= 12'h72f;
      20'h0d899: out <= 12'hfff;
      20'h0d89a: out <= 12'hfff;
      20'h0d89b: out <= 12'hc7f;
      20'h0d89c: out <= 12'h72f;
      20'h0d89d: out <= 12'hfff;
      20'h0d89e: out <= 12'hc7f;
      20'h0d89f: out <= 12'h000;
      20'h0d8a0: out <= 12'h000;
      20'h0d8a1: out <= 12'hbbb;
      20'h0d8a2: out <= 12'hfff;
      20'h0d8a3: out <= 12'hfff;
      20'h0d8a4: out <= 12'h666;
      20'h0d8a5: out <= 12'hfff;
      20'h0d8a6: out <= 12'hfff;
      20'h0d8a7: out <= 12'hfff;
      20'h0d8a8: out <= 12'hbbb;
      20'h0d8a9: out <= 12'hbbb;
      20'h0d8aa: out <= 12'h666;
      20'h0d8ab: out <= 12'h666;
      20'h0d8ac: out <= 12'hfff;
      20'h0d8ad: out <= 12'hfff;
      20'h0d8ae: out <= 12'hbbb;
      20'h0d8af: out <= 12'h000;
      20'h0d8b0: out <= 12'h000;
      20'h0d8b1: out <= 12'hbb0;
      20'h0d8b2: out <= 12'hee9;
      20'h0d8b3: out <= 12'hbb0;
      20'h0d8b4: out <= 12'hbb0;
      20'h0d8b5: out <= 12'h660;
      20'h0d8b6: out <= 12'h660;
      20'h0d8b7: out <= 12'h660;
      20'h0d8b8: out <= 12'hbb0;
      20'h0d8b9: out <= 12'h660;
      20'h0d8ba: out <= 12'h660;
      20'h0d8bb: out <= 12'hbb0;
      20'h0d8bc: out <= 12'hbb0;
      20'h0d8bd: out <= 12'hee9;
      20'h0d8be: out <= 12'hbb0;
      20'h0d8bf: out <= 12'h000;
      20'h0d8c0: out <= 12'h000;
      20'h0d8c1: out <= 12'h6af;
      20'h0d8c2: out <= 12'hfff;
      20'h0d8c3: out <= 12'hfff;
      20'h0d8c4: out <= 12'h6af;
      20'h0d8c5: out <= 12'h16d;
      20'h0d8c6: out <= 12'h16d;
      20'h0d8c7: out <= 12'hfff;
      20'h0d8c8: out <= 12'hfff;
      20'h0d8c9: out <= 12'h6af;
      20'h0d8ca: out <= 12'h16d;
      20'h0d8cb: out <= 12'h16d;
      20'h0d8cc: out <= 12'hfff;
      20'h0d8cd: out <= 12'hfff;
      20'h0d8ce: out <= 12'h6af;
      20'h0d8cf: out <= 12'h000;
      20'h0d8d0: out <= 12'h000;
      20'h0d8d1: out <= 12'hc7f;
      20'h0d8d2: out <= 12'hfff;
      20'h0d8d3: out <= 12'hc7f;
      20'h0d8d4: out <= 12'h72f;
      20'h0d8d5: out <= 12'hfff;
      20'h0d8d6: out <= 12'hfff;
      20'h0d8d7: out <= 12'hfff;
      20'h0d8d8: out <= 12'hfff;
      20'h0d8d9: out <= 12'hfff;
      20'h0d8da: out <= 12'hfff;
      20'h0d8db: out <= 12'h72f;
      20'h0d8dc: out <= 12'hc7f;
      20'h0d8dd: out <= 12'hfff;
      20'h0d8de: out <= 12'hc7f;
      20'h0d8df: out <= 12'h000;
      20'h0d8e0: out <= 12'h000;
      20'h0d8e1: out <= 12'hbbb;
      20'h0d8e2: out <= 12'hfff;
      20'h0d8e3: out <= 12'hfff;
      20'h0d8e4: out <= 12'hfff;
      20'h0d8e5: out <= 12'h666;
      20'h0d8e6: out <= 12'hbbb;
      20'h0d8e7: out <= 12'h666;
      20'h0d8e8: out <= 12'hbbb;
      20'h0d8e9: out <= 12'hbbb;
      20'h0d8ea: out <= 12'hfff;
      20'h0d8eb: out <= 12'hfff;
      20'h0d8ec: out <= 12'hfff;
      20'h0d8ed: out <= 12'hfff;
      20'h0d8ee: out <= 12'hbbb;
      20'h0d8ef: out <= 12'h000;
      20'h0d8f0: out <= 12'h000;
      20'h0d8f1: out <= 12'h6af;
      20'h0d8f2: out <= 12'hfff;
      20'h0d8f3: out <= 12'hfff;
      20'h0d8f4: out <= 12'hfff;
      20'h0d8f5: out <= 12'h6af;
      20'h0d8f6: out <= 12'h6af;
      20'h0d8f7: out <= 12'h16d;
      20'h0d8f8: out <= 12'h6af;
      20'h0d8f9: out <= 12'h16d;
      20'h0d8fa: out <= 12'h16d;
      20'h0d8fb: out <= 12'hfff;
      20'h0d8fc: out <= 12'hfff;
      20'h0d8fd: out <= 12'hfff;
      20'h0d8fe: out <= 12'h6af;
      20'h0d8ff: out <= 12'h000;
      20'h0d900: out <= 12'h000;
      20'h0d901: out <= 12'hbb0;
      20'h0d902: out <= 12'hee9;
      20'h0d903: out <= 12'hee9;
      20'h0d904: out <= 12'h660;
      20'h0d905: out <= 12'hbb0;
      20'h0d906: out <= 12'hee9;
      20'h0d907: out <= 12'hee9;
      20'h0d908: out <= 12'hee9;
      20'h0d909: out <= 12'hee9;
      20'h0d90a: out <= 12'hbb0;
      20'h0d90b: out <= 12'h660;
      20'h0d90c: out <= 12'hee9;
      20'h0d90d: out <= 12'hee9;
      20'h0d90e: out <= 12'hbb0;
      20'h0d90f: out <= 12'h000;
      20'h0d910: out <= 12'h603;
      20'h0d911: out <= 12'h603;
      20'h0d912: out <= 12'h603;
      20'h0d913: out <= 12'h603;
      20'h0d914: out <= 12'h603;
      20'h0d915: out <= 12'h603;
      20'h0d916: out <= 12'h603;
      20'h0d917: out <= 12'h603;
      20'h0d918: out <= 12'h603;
      20'h0d919: out <= 12'h603;
      20'h0d91a: out <= 12'h603;
      20'h0d91b: out <= 12'h603;
      20'h0d91c: out <= 12'h603;
      20'h0d91d: out <= 12'h603;
      20'h0d91e: out <= 12'h603;
      20'h0d91f: out <= 12'h603;
      20'h0d920: out <= 12'h603;
      20'h0d921: out <= 12'h603;
      20'h0d922: out <= 12'h603;
      20'h0d923: out <= 12'h603;
      20'h0d924: out <= 12'h603;
      20'h0d925: out <= 12'h603;
      20'h0d926: out <= 12'h603;
      20'h0d927: out <= 12'h603;
      20'h0d928: out <= 12'h603;
      20'h0d929: out <= 12'h603;
      20'h0d92a: out <= 12'h603;
      20'h0d92b: out <= 12'h603;
      20'h0d92c: out <= 12'h603;
      20'h0d92d: out <= 12'h603;
      20'h0d92e: out <= 12'h603;
      20'h0d92f: out <= 12'h603;
      20'h0d930: out <= 12'h603;
      20'h0d931: out <= 12'h603;
      20'h0d932: out <= 12'h603;
      20'h0d933: out <= 12'h603;
      20'h0d934: out <= 12'h603;
      20'h0d935: out <= 12'h603;
      20'h0d936: out <= 12'h603;
      20'h0d937: out <= 12'h603;
      20'h0d938: out <= 12'h603;
      20'h0d939: out <= 12'h603;
      20'h0d93a: out <= 12'h603;
      20'h0d93b: out <= 12'h603;
      20'h0d93c: out <= 12'h603;
      20'h0d93d: out <= 12'h603;
      20'h0d93e: out <= 12'h603;
      20'h0d93f: out <= 12'h603;
      20'h0d940: out <= 12'h603;
      20'h0d941: out <= 12'h603;
      20'h0d942: out <= 12'h603;
      20'h0d943: out <= 12'h603;
      20'h0d944: out <= 12'h603;
      20'h0d945: out <= 12'h603;
      20'h0d946: out <= 12'h603;
      20'h0d947: out <= 12'h603;
      20'h0d948: out <= 12'h603;
      20'h0d949: out <= 12'h603;
      20'h0d94a: out <= 12'h603;
      20'h0d94b: out <= 12'h603;
      20'h0d94c: out <= 12'h603;
      20'h0d94d: out <= 12'h603;
      20'h0d94e: out <= 12'h603;
      20'h0d94f: out <= 12'h603;
      20'h0d950: out <= 12'h603;
      20'h0d951: out <= 12'h603;
      20'h0d952: out <= 12'h603;
      20'h0d953: out <= 12'h603;
      20'h0d954: out <= 12'h603;
      20'h0d955: out <= 12'h603;
      20'h0d956: out <= 12'h603;
      20'h0d957: out <= 12'h603;
      20'h0d958: out <= 12'h603;
      20'h0d959: out <= 12'h603;
      20'h0d95a: out <= 12'h603;
      20'h0d95b: out <= 12'h603;
      20'h0d95c: out <= 12'h603;
      20'h0d95d: out <= 12'h603;
      20'h0d95e: out <= 12'h603;
      20'h0d95f: out <= 12'h603;
      20'h0d960: out <= 12'h603;
      20'h0d961: out <= 12'h603;
      20'h0d962: out <= 12'h603;
      20'h0d963: out <= 12'h603;
      20'h0d964: out <= 12'h603;
      20'h0d965: out <= 12'h603;
      20'h0d966: out <= 12'h603;
      20'h0d967: out <= 12'h603;
      20'h0d968: out <= 12'hee9;
      20'h0d969: out <= 12'hf87;
      20'h0d96a: out <= 12'hf87;
      20'h0d96b: out <= 12'hf87;
      20'h0d96c: out <= 12'hf87;
      20'h0d96d: out <= 12'hf87;
      20'h0d96e: out <= 12'hf87;
      20'h0d96f: out <= 12'hb27;
      20'h0d970: out <= 12'h000;
      20'h0d971: out <= 12'h000;
      20'h0d972: out <= 12'h000;
      20'h0d973: out <= 12'h000;
      20'h0d974: out <= 12'h000;
      20'h0d975: out <= 12'h000;
      20'h0d976: out <= 12'h000;
      20'h0d977: out <= 12'h000;
      20'h0d978: out <= 12'hbbb;
      20'h0d979: out <= 12'hbbb;
      20'h0d97a: out <= 12'hbbb;
      20'h0d97b: out <= 12'hbbb;
      20'h0d97c: out <= 12'hbbb;
      20'h0d97d: out <= 12'h000;
      20'h0d97e: out <= 12'hbbb;
      20'h0d97f: out <= 12'hbbb;
      20'h0d980: out <= 12'h000;
      20'h0d981: out <= 12'h000;
      20'h0d982: out <= 12'hbbb;
      20'h0d983: out <= 12'hbbb;
      20'h0d984: out <= 12'h000;
      20'h0d985: out <= 12'hbbb;
      20'h0d986: out <= 12'hbbb;
      20'h0d987: out <= 12'hbbb;
      20'h0d988: out <= 12'hbbb;
      20'h0d989: out <= 12'hbbb;
      20'h0d98a: out <= 12'h000;
      20'h0d98b: out <= 12'hbbb;
      20'h0d98c: out <= 12'hbbb;
      20'h0d98d: out <= 12'h000;
      20'h0d98e: out <= 12'hbbb;
      20'h0d98f: out <= 12'hbbb;
      20'h0d990: out <= 12'h000;
      20'h0d991: out <= 12'hbbb;
      20'h0d992: out <= 12'hbbb;
      20'h0d993: out <= 12'h000;
      20'h0d994: out <= 12'h000;
      20'h0d995: out <= 12'h000;
      20'h0d996: out <= 12'hbbb;
      20'h0d997: out <= 12'hbbb;
      20'h0d998: out <= 12'hbbb;
      20'h0d999: out <= 12'h000;
      20'h0d99a: out <= 12'h000;
      20'h0d99b: out <= 12'h000;
      20'h0d99c: out <= 12'h000;
      20'h0d99d: out <= 12'h000;
      20'h0d99e: out <= 12'h000;
      20'h0d99f: out <= 12'h000;
      20'h0d9a0: out <= 12'h000;
      20'h0d9a1: out <= 12'h000;
      20'h0d9a2: out <= 12'h000;
      20'h0d9a3: out <= 12'h000;
      20'h0d9a4: out <= 12'h000;
      20'h0d9a5: out <= 12'h000;
      20'h0d9a6: out <= 12'h000;
      20'h0d9a7: out <= 12'h000;
      20'h0d9a8: out <= 12'h000;
      20'h0d9a9: out <= 12'hc7f;
      20'h0d9aa: out <= 12'hfff;
      20'h0d9ab: out <= 12'h72f;
      20'h0d9ac: out <= 12'hc7f;
      20'h0d9ad: out <= 12'hfff;
      20'h0d9ae: out <= 12'hfff;
      20'h0d9af: out <= 12'hfff;
      20'h0d9b0: out <= 12'h72f;
      20'h0d9b1: out <= 12'hfff;
      20'h0d9b2: out <= 12'hfff;
      20'h0d9b3: out <= 12'hc7f;
      20'h0d9b4: out <= 12'h72f;
      20'h0d9b5: out <= 12'hfff;
      20'h0d9b6: out <= 12'hc7f;
      20'h0d9b7: out <= 12'h000;
      20'h0d9b8: out <= 12'h000;
      20'h0d9b9: out <= 12'hbbb;
      20'h0d9ba: out <= 12'hfff;
      20'h0d9bb: out <= 12'h666;
      20'h0d9bc: out <= 12'hfff;
      20'h0d9bd: out <= 12'hfff;
      20'h0d9be: out <= 12'hbbb;
      20'h0d9bf: out <= 12'hbbb;
      20'h0d9c0: out <= 12'hbbb;
      20'h0d9c1: out <= 12'hbbb;
      20'h0d9c2: out <= 12'hbbb;
      20'h0d9c3: out <= 12'h666;
      20'h0d9c4: out <= 12'h666;
      20'h0d9c5: out <= 12'hfff;
      20'h0d9c6: out <= 12'hbbb;
      20'h0d9c7: out <= 12'h000;
      20'h0d9c8: out <= 12'h000;
      20'h0d9c9: out <= 12'hbb0;
      20'h0d9ca: out <= 12'hee9;
      20'h0d9cb: out <= 12'h660;
      20'h0d9cc: out <= 12'h660;
      20'h0d9cd: out <= 12'h660;
      20'h0d9ce: out <= 12'h660;
      20'h0d9cf: out <= 12'h660;
      20'h0d9d0: out <= 12'hbb0;
      20'h0d9d1: out <= 12'h660;
      20'h0d9d2: out <= 12'h660;
      20'h0d9d3: out <= 12'h660;
      20'h0d9d4: out <= 12'h660;
      20'h0d9d5: out <= 12'hee9;
      20'h0d9d6: out <= 12'hbb0;
      20'h0d9d7: out <= 12'h000;
      20'h0d9d8: out <= 12'h000;
      20'h0d9d9: out <= 12'h6af;
      20'h0d9da: out <= 12'hfff;
      20'h0d9db: out <= 12'hfff;
      20'h0d9dc: out <= 12'h6af;
      20'h0d9dd: out <= 12'h16d;
      20'h0d9de: out <= 12'h16d;
      20'h0d9df: out <= 12'hfff;
      20'h0d9e0: out <= 12'hfff;
      20'h0d9e1: out <= 12'h6af;
      20'h0d9e2: out <= 12'h16d;
      20'h0d9e3: out <= 12'h16d;
      20'h0d9e4: out <= 12'hfff;
      20'h0d9e5: out <= 12'hfff;
      20'h0d9e6: out <= 12'h6af;
      20'h0d9e7: out <= 12'h000;
      20'h0d9e8: out <= 12'h000;
      20'h0d9e9: out <= 12'hc7f;
      20'h0d9ea: out <= 12'hfff;
      20'h0d9eb: out <= 12'hc7f;
      20'h0d9ec: out <= 12'h72f;
      20'h0d9ed: out <= 12'hc7f;
      20'h0d9ee: out <= 12'hc7f;
      20'h0d9ef: out <= 12'hc7f;
      20'h0d9f0: out <= 12'hc7f;
      20'h0d9f1: out <= 12'hc7f;
      20'h0d9f2: out <= 12'hc7f;
      20'h0d9f3: out <= 12'h72f;
      20'h0d9f4: out <= 12'hc7f;
      20'h0d9f5: out <= 12'hfff;
      20'h0d9f6: out <= 12'hc7f;
      20'h0d9f7: out <= 12'h000;
      20'h0d9f8: out <= 12'h000;
      20'h0d9f9: out <= 12'hbbb;
      20'h0d9fa: out <= 12'hfff;
      20'h0d9fb: out <= 12'hfff;
      20'h0d9fc: out <= 12'hfff;
      20'h0d9fd: out <= 12'h666;
      20'h0d9fe: out <= 12'hbbb;
      20'h0d9ff: out <= 12'h666;
      20'h0da00: out <= 12'h666;
      20'h0da01: out <= 12'hbbb;
      20'h0da02: out <= 12'hbbb;
      20'h0da03: out <= 12'hfff;
      20'h0da04: out <= 12'hfff;
      20'h0da05: out <= 12'hfff;
      20'h0da06: out <= 12'hbbb;
      20'h0da07: out <= 12'h000;
      20'h0da08: out <= 12'h000;
      20'h0da09: out <= 12'h6af;
      20'h0da0a: out <= 12'hfff;
      20'h0da0b: out <= 12'hfff;
      20'h0da0c: out <= 12'hfff;
      20'h0da0d: out <= 12'h6af;
      20'h0da0e: out <= 12'h6af;
      20'h0da0f: out <= 12'h16d;
      20'h0da10: out <= 12'h6af;
      20'h0da11: out <= 12'h16d;
      20'h0da12: out <= 12'h16d;
      20'h0da13: out <= 12'hfff;
      20'h0da14: out <= 12'hfff;
      20'h0da15: out <= 12'hfff;
      20'h0da16: out <= 12'h6af;
      20'h0da17: out <= 12'h000;
      20'h0da18: out <= 12'h000;
      20'h0da19: out <= 12'hbb0;
      20'h0da1a: out <= 12'hee9;
      20'h0da1b: out <= 12'hee9;
      20'h0da1c: out <= 12'h660;
      20'h0da1d: out <= 12'hbb0;
      20'h0da1e: out <= 12'hee9;
      20'h0da1f: out <= 12'hee9;
      20'h0da20: out <= 12'hee9;
      20'h0da21: out <= 12'hee9;
      20'h0da22: out <= 12'hbb0;
      20'h0da23: out <= 12'h660;
      20'h0da24: out <= 12'hee9;
      20'h0da25: out <= 12'hee9;
      20'h0da26: out <= 12'hbb0;
      20'h0da27: out <= 12'h000;
      20'h0da28: out <= 12'h603;
      20'h0da29: out <= 12'h603;
      20'h0da2a: out <= 12'h603;
      20'h0da2b: out <= 12'h603;
      20'h0da2c: out <= 12'h603;
      20'h0da2d: out <= 12'h603;
      20'h0da2e: out <= 12'h603;
      20'h0da2f: out <= 12'h603;
      20'h0da30: out <= 12'h603;
      20'h0da31: out <= 12'h603;
      20'h0da32: out <= 12'h603;
      20'h0da33: out <= 12'h603;
      20'h0da34: out <= 12'h603;
      20'h0da35: out <= 12'h603;
      20'h0da36: out <= 12'h603;
      20'h0da37: out <= 12'h603;
      20'h0da38: out <= 12'h603;
      20'h0da39: out <= 12'h603;
      20'h0da3a: out <= 12'h603;
      20'h0da3b: out <= 12'h603;
      20'h0da3c: out <= 12'h603;
      20'h0da3d: out <= 12'h603;
      20'h0da3e: out <= 12'h603;
      20'h0da3f: out <= 12'h603;
      20'h0da40: out <= 12'h603;
      20'h0da41: out <= 12'h603;
      20'h0da42: out <= 12'h603;
      20'h0da43: out <= 12'h603;
      20'h0da44: out <= 12'h603;
      20'h0da45: out <= 12'h603;
      20'h0da46: out <= 12'h603;
      20'h0da47: out <= 12'h603;
      20'h0da48: out <= 12'h603;
      20'h0da49: out <= 12'h603;
      20'h0da4a: out <= 12'h603;
      20'h0da4b: out <= 12'h603;
      20'h0da4c: out <= 12'h603;
      20'h0da4d: out <= 12'h603;
      20'h0da4e: out <= 12'h603;
      20'h0da4f: out <= 12'h603;
      20'h0da50: out <= 12'h603;
      20'h0da51: out <= 12'h603;
      20'h0da52: out <= 12'h603;
      20'h0da53: out <= 12'h603;
      20'h0da54: out <= 12'h603;
      20'h0da55: out <= 12'h603;
      20'h0da56: out <= 12'h603;
      20'h0da57: out <= 12'h603;
      20'h0da58: out <= 12'h603;
      20'h0da59: out <= 12'h603;
      20'h0da5a: out <= 12'h603;
      20'h0da5b: out <= 12'h603;
      20'h0da5c: out <= 12'h603;
      20'h0da5d: out <= 12'h603;
      20'h0da5e: out <= 12'h603;
      20'h0da5f: out <= 12'h603;
      20'h0da60: out <= 12'h603;
      20'h0da61: out <= 12'h603;
      20'h0da62: out <= 12'h603;
      20'h0da63: out <= 12'h603;
      20'h0da64: out <= 12'h603;
      20'h0da65: out <= 12'h603;
      20'h0da66: out <= 12'h603;
      20'h0da67: out <= 12'h603;
      20'h0da68: out <= 12'h603;
      20'h0da69: out <= 12'h603;
      20'h0da6a: out <= 12'h603;
      20'h0da6b: out <= 12'h603;
      20'h0da6c: out <= 12'h603;
      20'h0da6d: out <= 12'h603;
      20'h0da6e: out <= 12'h603;
      20'h0da6f: out <= 12'h603;
      20'h0da70: out <= 12'h603;
      20'h0da71: out <= 12'h603;
      20'h0da72: out <= 12'h603;
      20'h0da73: out <= 12'h603;
      20'h0da74: out <= 12'h603;
      20'h0da75: out <= 12'h603;
      20'h0da76: out <= 12'h603;
      20'h0da77: out <= 12'h603;
      20'h0da78: out <= 12'h603;
      20'h0da79: out <= 12'h603;
      20'h0da7a: out <= 12'h603;
      20'h0da7b: out <= 12'h603;
      20'h0da7c: out <= 12'h603;
      20'h0da7d: out <= 12'h603;
      20'h0da7e: out <= 12'h603;
      20'h0da7f: out <= 12'h603;
      20'h0da80: out <= 12'hb27;
      20'h0da81: out <= 12'hb27;
      20'h0da82: out <= 12'hb27;
      20'h0da83: out <= 12'hb27;
      20'h0da84: out <= 12'hb27;
      20'h0da85: out <= 12'hb27;
      20'h0da86: out <= 12'hb27;
      20'h0da87: out <= 12'hb27;
      20'h0da88: out <= 12'h000;
      20'h0da89: out <= 12'h000;
      20'h0da8a: out <= 12'h000;
      20'h0da8b: out <= 12'h000;
      20'h0da8c: out <= 12'h000;
      20'h0da8d: out <= 12'h000;
      20'h0da8e: out <= 12'h000;
      20'h0da8f: out <= 12'h000;
      20'h0da90: out <= 12'h000;
      20'h0da91: out <= 12'h000;
      20'h0da92: out <= 12'h000;
      20'h0da93: out <= 12'h000;
      20'h0da94: out <= 12'h000;
      20'h0da95: out <= 12'h000;
      20'h0da96: out <= 12'h000;
      20'h0da97: out <= 12'h000;
      20'h0da98: out <= 12'h000;
      20'h0da99: out <= 12'h000;
      20'h0da9a: out <= 12'h000;
      20'h0da9b: out <= 12'h000;
      20'h0da9c: out <= 12'h000;
      20'h0da9d: out <= 12'h000;
      20'h0da9e: out <= 12'h000;
      20'h0da9f: out <= 12'h000;
      20'h0daa0: out <= 12'h000;
      20'h0daa1: out <= 12'h000;
      20'h0daa2: out <= 12'h000;
      20'h0daa3: out <= 12'h000;
      20'h0daa4: out <= 12'h000;
      20'h0daa5: out <= 12'h000;
      20'h0daa6: out <= 12'h000;
      20'h0daa7: out <= 12'h000;
      20'h0daa8: out <= 12'h000;
      20'h0daa9: out <= 12'h000;
      20'h0daaa: out <= 12'h000;
      20'h0daab: out <= 12'h000;
      20'h0daac: out <= 12'h000;
      20'h0daad: out <= 12'h000;
      20'h0daae: out <= 12'h000;
      20'h0daaf: out <= 12'h000;
      20'h0dab0: out <= 12'h000;
      20'h0dab1: out <= 12'h000;
      20'h0dab2: out <= 12'h000;
      20'h0dab3: out <= 12'h000;
      20'h0dab4: out <= 12'h000;
      20'h0dab5: out <= 12'h000;
      20'h0dab6: out <= 12'h000;
      20'h0dab7: out <= 12'h000;
      20'h0dab8: out <= 12'h000;
      20'h0dab9: out <= 12'h000;
      20'h0daba: out <= 12'h000;
      20'h0dabb: out <= 12'h000;
      20'h0dabc: out <= 12'h000;
      20'h0dabd: out <= 12'h000;
      20'h0dabe: out <= 12'h000;
      20'h0dabf: out <= 12'h000;
      20'h0dac0: out <= 12'h000;
      20'h0dac1: out <= 12'hc7f;
      20'h0dac2: out <= 12'hfff;
      20'h0dac3: out <= 12'h72f;
      20'h0dac4: out <= 12'hc7f;
      20'h0dac5: out <= 12'h72f;
      20'h0dac6: out <= 12'h72f;
      20'h0dac7: out <= 12'h72f;
      20'h0dac8: out <= 12'h72f;
      20'h0dac9: out <= 12'hfff;
      20'h0daca: out <= 12'hfff;
      20'h0dacb: out <= 12'hc7f;
      20'h0dacc: out <= 12'h72f;
      20'h0dacd: out <= 12'hfff;
      20'h0dace: out <= 12'hc7f;
      20'h0dacf: out <= 12'h000;
      20'h0dad0: out <= 12'h000;
      20'h0dad1: out <= 12'hbbb;
      20'h0dad2: out <= 12'hfff;
      20'h0dad3: out <= 12'h666;
      20'h0dad4: out <= 12'hfff;
      20'h0dad5: out <= 12'hbbb;
      20'h0dad6: out <= 12'hbbb;
      20'h0dad7: out <= 12'hbbb;
      20'h0dad8: out <= 12'hbbb;
      20'h0dad9: out <= 12'h666;
      20'h0dada: out <= 12'h666;
      20'h0dadb: out <= 12'h666;
      20'h0dadc: out <= 12'h666;
      20'h0dadd: out <= 12'hfff;
      20'h0dade: out <= 12'hbbb;
      20'h0dadf: out <= 12'h000;
      20'h0dae0: out <= 12'h000;
      20'h0dae1: out <= 12'hbb0;
      20'h0dae2: out <= 12'hee9;
      20'h0dae3: out <= 12'hbb0;
      20'h0dae4: out <= 12'hbb0;
      20'h0dae5: out <= 12'h660;
      20'h0dae6: out <= 12'hbb0;
      20'h0dae7: out <= 12'hee9;
      20'h0dae8: out <= 12'hee9;
      20'h0dae9: out <= 12'hbb0;
      20'h0daea: out <= 12'h660;
      20'h0daeb: out <= 12'hbb0;
      20'h0daec: out <= 12'hbb0;
      20'h0daed: out <= 12'hee9;
      20'h0daee: out <= 12'hbb0;
      20'h0daef: out <= 12'h000;
      20'h0daf0: out <= 12'h000;
      20'h0daf1: out <= 12'h6af;
      20'h0daf2: out <= 12'hfff;
      20'h0daf3: out <= 12'hfff;
      20'h0daf4: out <= 12'h6af;
      20'h0daf5: out <= 12'h16d;
      20'h0daf6: out <= 12'h16d;
      20'h0daf7: out <= 12'hfff;
      20'h0daf8: out <= 12'hfff;
      20'h0daf9: out <= 12'h6af;
      20'h0dafa: out <= 12'h16d;
      20'h0dafb: out <= 12'h16d;
      20'h0dafc: out <= 12'hfff;
      20'h0dafd: out <= 12'hfff;
      20'h0dafe: out <= 12'h6af;
      20'h0daff: out <= 12'h000;
      20'h0db00: out <= 12'h000;
      20'h0db01: out <= 12'hc7f;
      20'h0db02: out <= 12'hfff;
      20'h0db03: out <= 12'hc7f;
      20'h0db04: out <= 12'h72f;
      20'h0db05: out <= 12'h72f;
      20'h0db06: out <= 12'h72f;
      20'h0db07: out <= 12'h72f;
      20'h0db08: out <= 12'h72f;
      20'h0db09: out <= 12'h72f;
      20'h0db0a: out <= 12'h72f;
      20'h0db0b: out <= 12'h72f;
      20'h0db0c: out <= 12'hc7f;
      20'h0db0d: out <= 12'hfff;
      20'h0db0e: out <= 12'hc7f;
      20'h0db0f: out <= 12'h000;
      20'h0db10: out <= 12'h000;
      20'h0db11: out <= 12'hbbb;
      20'h0db12: out <= 12'hfff;
      20'h0db13: out <= 12'hfff;
      20'h0db14: out <= 12'hfff;
      20'h0db15: out <= 12'h666;
      20'h0db16: out <= 12'hbbb;
      20'h0db17: out <= 12'h666;
      20'h0db18: out <= 12'h666;
      20'h0db19: out <= 12'h666;
      20'h0db1a: out <= 12'hbbb;
      20'h0db1b: out <= 12'hbbb;
      20'h0db1c: out <= 12'hfff;
      20'h0db1d: out <= 12'hfff;
      20'h0db1e: out <= 12'hbbb;
      20'h0db1f: out <= 12'h000;
      20'h0db20: out <= 12'h000;
      20'h0db21: out <= 12'h6af;
      20'h0db22: out <= 12'hfff;
      20'h0db23: out <= 12'hfff;
      20'h0db24: out <= 12'hfff;
      20'h0db25: out <= 12'h6af;
      20'h0db26: out <= 12'h6af;
      20'h0db27: out <= 12'h16d;
      20'h0db28: out <= 12'h6af;
      20'h0db29: out <= 12'h16d;
      20'h0db2a: out <= 12'h16d;
      20'h0db2b: out <= 12'hfff;
      20'h0db2c: out <= 12'hfff;
      20'h0db2d: out <= 12'hfff;
      20'h0db2e: out <= 12'h6af;
      20'h0db2f: out <= 12'h000;
      20'h0db30: out <= 12'h000;
      20'h0db31: out <= 12'hbb0;
      20'h0db32: out <= 12'hee9;
      20'h0db33: out <= 12'hee9;
      20'h0db34: out <= 12'h660;
      20'h0db35: out <= 12'hbb0;
      20'h0db36: out <= 12'hbb0;
      20'h0db37: out <= 12'hee9;
      20'h0db38: out <= 12'hee9;
      20'h0db39: out <= 12'hbb0;
      20'h0db3a: out <= 12'hbb0;
      20'h0db3b: out <= 12'h660;
      20'h0db3c: out <= 12'hee9;
      20'h0db3d: out <= 12'hee9;
      20'h0db3e: out <= 12'hbb0;
      20'h0db3f: out <= 12'h000;
      20'h0db40: out <= 12'h603;
      20'h0db41: out <= 12'h603;
      20'h0db42: out <= 12'h603;
      20'h0db43: out <= 12'h603;
      20'h0db44: out <= 12'h603;
      20'h0db45: out <= 12'h603;
      20'h0db46: out <= 12'h603;
      20'h0db47: out <= 12'h603;
      20'h0db48: out <= 12'h603;
      20'h0db49: out <= 12'h603;
      20'h0db4a: out <= 12'h603;
      20'h0db4b: out <= 12'h603;
      20'h0db4c: out <= 12'h603;
      20'h0db4d: out <= 12'h603;
      20'h0db4e: out <= 12'h603;
      20'h0db4f: out <= 12'h603;
      20'h0db50: out <= 12'h603;
      20'h0db51: out <= 12'h603;
      20'h0db52: out <= 12'h603;
      20'h0db53: out <= 12'h603;
      20'h0db54: out <= 12'h603;
      20'h0db55: out <= 12'h603;
      20'h0db56: out <= 12'h603;
      20'h0db57: out <= 12'h603;
      20'h0db58: out <= 12'h603;
      20'h0db59: out <= 12'h603;
      20'h0db5a: out <= 12'h603;
      20'h0db5b: out <= 12'h603;
      20'h0db5c: out <= 12'h603;
      20'h0db5d: out <= 12'h603;
      20'h0db5e: out <= 12'h603;
      20'h0db5f: out <= 12'h603;
      20'h0db60: out <= 12'h603;
      20'h0db61: out <= 12'h603;
      20'h0db62: out <= 12'h603;
      20'h0db63: out <= 12'h603;
      20'h0db64: out <= 12'h603;
      20'h0db65: out <= 12'h603;
      20'h0db66: out <= 12'h603;
      20'h0db67: out <= 12'h603;
      20'h0db68: out <= 12'h603;
      20'h0db69: out <= 12'h603;
      20'h0db6a: out <= 12'h603;
      20'h0db6b: out <= 12'h603;
      20'h0db6c: out <= 12'h603;
      20'h0db6d: out <= 12'h603;
      20'h0db6e: out <= 12'h603;
      20'h0db6f: out <= 12'h603;
      20'h0db70: out <= 12'h603;
      20'h0db71: out <= 12'h603;
      20'h0db72: out <= 12'h603;
      20'h0db73: out <= 12'h603;
      20'h0db74: out <= 12'h603;
      20'h0db75: out <= 12'h603;
      20'h0db76: out <= 12'h603;
      20'h0db77: out <= 12'h603;
      20'h0db78: out <= 12'h603;
      20'h0db79: out <= 12'h603;
      20'h0db7a: out <= 12'h603;
      20'h0db7b: out <= 12'h603;
      20'h0db7c: out <= 12'h603;
      20'h0db7d: out <= 12'h603;
      20'h0db7e: out <= 12'h603;
      20'h0db7f: out <= 12'h603;
      20'h0db80: out <= 12'h603;
      20'h0db81: out <= 12'h603;
      20'h0db82: out <= 12'h603;
      20'h0db83: out <= 12'h603;
      20'h0db84: out <= 12'h603;
      20'h0db85: out <= 12'h603;
      20'h0db86: out <= 12'h603;
      20'h0db87: out <= 12'h603;
      20'h0db88: out <= 12'h603;
      20'h0db89: out <= 12'h603;
      20'h0db8a: out <= 12'h603;
      20'h0db8b: out <= 12'h603;
      20'h0db8c: out <= 12'h603;
      20'h0db8d: out <= 12'h603;
      20'h0db8e: out <= 12'h603;
      20'h0db8f: out <= 12'h603;
      20'h0db90: out <= 12'h603;
      20'h0db91: out <= 12'h603;
      20'h0db92: out <= 12'h603;
      20'h0db93: out <= 12'h603;
      20'h0db94: out <= 12'h603;
      20'h0db95: out <= 12'h603;
      20'h0db96: out <= 12'h603;
      20'h0db97: out <= 12'h603;
      20'h0db98: out <= 12'hee9;
      20'h0db99: out <= 12'hee9;
      20'h0db9a: out <= 12'hee9;
      20'h0db9b: out <= 12'hee9;
      20'h0db9c: out <= 12'hee9;
      20'h0db9d: out <= 12'hee9;
      20'h0db9e: out <= 12'hee9;
      20'h0db9f: out <= 12'hb27;
      20'h0dba0: out <= 12'h000;
      20'h0dba1: out <= 12'h000;
      20'h0dba2: out <= 12'h000;
      20'h0dba3: out <= 12'h000;
      20'h0dba4: out <= 12'h000;
      20'h0dba5: out <= 12'h000;
      20'h0dba6: out <= 12'h000;
      20'h0dba7: out <= 12'h000;
      20'h0dba8: out <= 12'h000;
      20'h0dba9: out <= 12'h000;
      20'h0dbaa: out <= 12'h000;
      20'h0dbab: out <= 12'h000;
      20'h0dbac: out <= 12'h000;
      20'h0dbad: out <= 12'h000;
      20'h0dbae: out <= 12'h666;
      20'h0dbaf: out <= 12'hbbb;
      20'h0dbb0: out <= 12'hfff;
      20'h0dbb1: out <= 12'hbbb;
      20'h0dbb2: out <= 12'h666;
      20'h0dbb3: out <= 12'h000;
      20'h0dbb4: out <= 12'h000;
      20'h0dbb5: out <= 12'h000;
      20'h0dbb6: out <= 12'h000;
      20'h0dbb7: out <= 12'h000;
      20'h0dbb8: out <= 12'h000;
      20'h0dbb9: out <= 12'h000;
      20'h0dbba: out <= 12'h000;
      20'h0dbbb: out <= 12'h000;
      20'h0dbbc: out <= 12'h000;
      20'h0dbbd: out <= 12'h000;
      20'h0dbbe: out <= 12'h000;
      20'h0dbbf: out <= 12'h000;
      20'h0dbc0: out <= 12'h000;
      20'h0dbc1: out <= 12'h000;
      20'h0dbc2: out <= 12'h000;
      20'h0dbc3: out <= 12'h000;
      20'h0dbc4: out <= 12'h000;
      20'h0dbc5: out <= 12'h000;
      20'h0dbc6: out <= 12'h000;
      20'h0dbc7: out <= 12'h000;
      20'h0dbc8: out <= 12'h000;
      20'h0dbc9: out <= 12'h000;
      20'h0dbca: out <= 12'h000;
      20'h0dbcb: out <= 12'h000;
      20'h0dbcc: out <= 12'h000;
      20'h0dbcd: out <= 12'h000;
      20'h0dbce: out <= 12'h000;
      20'h0dbcf: out <= 12'h000;
      20'h0dbd0: out <= 12'h000;
      20'h0dbd1: out <= 12'h000;
      20'h0dbd2: out <= 12'h000;
      20'h0dbd3: out <= 12'h000;
      20'h0dbd4: out <= 12'h000;
      20'h0dbd5: out <= 12'h000;
      20'h0dbd6: out <= 12'h000;
      20'h0dbd7: out <= 12'h000;
      20'h0dbd8: out <= 12'h000;
      20'h0dbd9: out <= 12'hc7f;
      20'h0dbda: out <= 12'hfff;
      20'h0dbdb: out <= 12'h72f;
      20'h0dbdc: out <= 12'hc7f;
      20'h0dbdd: out <= 12'hfff;
      20'h0dbde: out <= 12'hfff;
      20'h0dbdf: out <= 12'hfff;
      20'h0dbe0: out <= 12'hfff;
      20'h0dbe1: out <= 12'hfff;
      20'h0dbe2: out <= 12'hfff;
      20'h0dbe3: out <= 12'hc7f;
      20'h0dbe4: out <= 12'h72f;
      20'h0dbe5: out <= 12'hfff;
      20'h0dbe6: out <= 12'hc7f;
      20'h0dbe7: out <= 12'h000;
      20'h0dbe8: out <= 12'h000;
      20'h0dbe9: out <= 12'hbbb;
      20'h0dbea: out <= 12'hfff;
      20'h0dbeb: out <= 12'h666;
      20'h0dbec: out <= 12'hfff;
      20'h0dbed: out <= 12'hbbb;
      20'h0dbee: out <= 12'hbbb;
      20'h0dbef: out <= 12'hbbb;
      20'h0dbf0: out <= 12'h666;
      20'h0dbf1: out <= 12'h666;
      20'h0dbf2: out <= 12'h666;
      20'h0dbf3: out <= 12'h666;
      20'h0dbf4: out <= 12'h666;
      20'h0dbf5: out <= 12'hfff;
      20'h0dbf6: out <= 12'hbbb;
      20'h0dbf7: out <= 12'h000;
      20'h0dbf8: out <= 12'h000;
      20'h0dbf9: out <= 12'hbb0;
      20'h0dbfa: out <= 12'hee9;
      20'h0dbfb: out <= 12'h660;
      20'h0dbfc: out <= 12'h660;
      20'h0dbfd: out <= 12'h660;
      20'h0dbfe: out <= 12'hbb0;
      20'h0dbff: out <= 12'hee9;
      20'h0dc00: out <= 12'hee9;
      20'h0dc01: out <= 12'hbb0;
      20'h0dc02: out <= 12'h660;
      20'h0dc03: out <= 12'h660;
      20'h0dc04: out <= 12'h660;
      20'h0dc05: out <= 12'hee9;
      20'h0dc06: out <= 12'hbb0;
      20'h0dc07: out <= 12'h000;
      20'h0dc08: out <= 12'h000;
      20'h0dc09: out <= 12'h6af;
      20'h0dc0a: out <= 12'hfff;
      20'h0dc0b: out <= 12'hfff;
      20'h0dc0c: out <= 12'h6af;
      20'h0dc0d: out <= 12'h16d;
      20'h0dc0e: out <= 12'h16d;
      20'h0dc0f: out <= 12'hfff;
      20'h0dc10: out <= 12'hfff;
      20'h0dc11: out <= 12'h6af;
      20'h0dc12: out <= 12'h16d;
      20'h0dc13: out <= 12'h16d;
      20'h0dc14: out <= 12'hfff;
      20'h0dc15: out <= 12'hfff;
      20'h0dc16: out <= 12'h6af;
      20'h0dc17: out <= 12'h000;
      20'h0dc18: out <= 12'h000;
      20'h0dc19: out <= 12'hc7f;
      20'h0dc1a: out <= 12'hfff;
      20'h0dc1b: out <= 12'hc7f;
      20'h0dc1c: out <= 12'h72f;
      20'h0dc1d: out <= 12'h72f;
      20'h0dc1e: out <= 12'h72f;
      20'h0dc1f: out <= 12'h72f;
      20'h0dc20: out <= 12'h72f;
      20'h0dc21: out <= 12'h72f;
      20'h0dc22: out <= 12'h72f;
      20'h0dc23: out <= 12'h72f;
      20'h0dc24: out <= 12'hc7f;
      20'h0dc25: out <= 12'hfff;
      20'h0dc26: out <= 12'hc7f;
      20'h0dc27: out <= 12'h000;
      20'h0dc28: out <= 12'h000;
      20'h0dc29: out <= 12'hbbb;
      20'h0dc2a: out <= 12'hfff;
      20'h0dc2b: out <= 12'hfff;
      20'h0dc2c: out <= 12'hfff;
      20'h0dc2d: out <= 12'h666;
      20'h0dc2e: out <= 12'hbbb;
      20'h0dc2f: out <= 12'hfff;
      20'h0dc30: out <= 12'hfff;
      20'h0dc31: out <= 12'hfff;
      20'h0dc32: out <= 12'hfff;
      20'h0dc33: out <= 12'hfff;
      20'h0dc34: out <= 12'hfff;
      20'h0dc35: out <= 12'hfff;
      20'h0dc36: out <= 12'hbbb;
      20'h0dc37: out <= 12'h000;
      20'h0dc38: out <= 12'h000;
      20'h0dc39: out <= 12'h6af;
      20'h0dc3a: out <= 12'hfff;
      20'h0dc3b: out <= 12'hfff;
      20'h0dc3c: out <= 12'hfff;
      20'h0dc3d: out <= 12'h6af;
      20'h0dc3e: out <= 12'h6af;
      20'h0dc3f: out <= 12'h16d;
      20'h0dc40: out <= 12'h6af;
      20'h0dc41: out <= 12'h16d;
      20'h0dc42: out <= 12'h16d;
      20'h0dc43: out <= 12'hfff;
      20'h0dc44: out <= 12'hfff;
      20'h0dc45: out <= 12'hfff;
      20'h0dc46: out <= 12'h6af;
      20'h0dc47: out <= 12'h000;
      20'h0dc48: out <= 12'h000;
      20'h0dc49: out <= 12'hbb0;
      20'h0dc4a: out <= 12'hee9;
      20'h0dc4b: out <= 12'hee9;
      20'h0dc4c: out <= 12'hee9;
      20'h0dc4d: out <= 12'h660;
      20'h0dc4e: out <= 12'hbb0;
      20'h0dc4f: out <= 12'hee9;
      20'h0dc50: out <= 12'hee9;
      20'h0dc51: out <= 12'hbb0;
      20'h0dc52: out <= 12'h660;
      20'h0dc53: out <= 12'hee9;
      20'h0dc54: out <= 12'hee9;
      20'h0dc55: out <= 12'hee9;
      20'h0dc56: out <= 12'hbb0;
      20'h0dc57: out <= 12'h000;
      20'h0dc58: out <= 12'h603;
      20'h0dc59: out <= 12'h603;
      20'h0dc5a: out <= 12'h603;
      20'h0dc5b: out <= 12'h603;
      20'h0dc5c: out <= 12'h603;
      20'h0dc5d: out <= 12'h603;
      20'h0dc5e: out <= 12'h603;
      20'h0dc5f: out <= 12'h603;
      20'h0dc60: out <= 12'h603;
      20'h0dc61: out <= 12'h603;
      20'h0dc62: out <= 12'h603;
      20'h0dc63: out <= 12'h603;
      20'h0dc64: out <= 12'h603;
      20'h0dc65: out <= 12'h603;
      20'h0dc66: out <= 12'h603;
      20'h0dc67: out <= 12'h603;
      20'h0dc68: out <= 12'h603;
      20'h0dc69: out <= 12'h603;
      20'h0dc6a: out <= 12'h603;
      20'h0dc6b: out <= 12'h603;
      20'h0dc6c: out <= 12'h603;
      20'h0dc6d: out <= 12'h603;
      20'h0dc6e: out <= 12'h603;
      20'h0dc6f: out <= 12'h603;
      20'h0dc70: out <= 12'h603;
      20'h0dc71: out <= 12'h603;
      20'h0dc72: out <= 12'h603;
      20'h0dc73: out <= 12'h603;
      20'h0dc74: out <= 12'h603;
      20'h0dc75: out <= 12'h603;
      20'h0dc76: out <= 12'h603;
      20'h0dc77: out <= 12'h603;
      20'h0dc78: out <= 12'h603;
      20'h0dc79: out <= 12'h603;
      20'h0dc7a: out <= 12'h603;
      20'h0dc7b: out <= 12'h603;
      20'h0dc7c: out <= 12'h603;
      20'h0dc7d: out <= 12'h603;
      20'h0dc7e: out <= 12'h603;
      20'h0dc7f: out <= 12'h603;
      20'h0dc80: out <= 12'h603;
      20'h0dc81: out <= 12'h603;
      20'h0dc82: out <= 12'h603;
      20'h0dc83: out <= 12'h603;
      20'h0dc84: out <= 12'h603;
      20'h0dc85: out <= 12'h603;
      20'h0dc86: out <= 12'h603;
      20'h0dc87: out <= 12'h603;
      20'h0dc88: out <= 12'h603;
      20'h0dc89: out <= 12'h603;
      20'h0dc8a: out <= 12'h603;
      20'h0dc8b: out <= 12'h603;
      20'h0dc8c: out <= 12'h603;
      20'h0dc8d: out <= 12'h603;
      20'h0dc8e: out <= 12'h603;
      20'h0dc8f: out <= 12'h603;
      20'h0dc90: out <= 12'h603;
      20'h0dc91: out <= 12'h603;
      20'h0dc92: out <= 12'h603;
      20'h0dc93: out <= 12'h603;
      20'h0dc94: out <= 12'h603;
      20'h0dc95: out <= 12'h603;
      20'h0dc96: out <= 12'h603;
      20'h0dc97: out <= 12'h603;
      20'h0dc98: out <= 12'h603;
      20'h0dc99: out <= 12'h603;
      20'h0dc9a: out <= 12'h603;
      20'h0dc9b: out <= 12'h603;
      20'h0dc9c: out <= 12'h603;
      20'h0dc9d: out <= 12'h603;
      20'h0dc9e: out <= 12'h603;
      20'h0dc9f: out <= 12'h603;
      20'h0dca0: out <= 12'h603;
      20'h0dca1: out <= 12'h603;
      20'h0dca2: out <= 12'h603;
      20'h0dca3: out <= 12'h603;
      20'h0dca4: out <= 12'h603;
      20'h0dca5: out <= 12'h603;
      20'h0dca6: out <= 12'h603;
      20'h0dca7: out <= 12'h603;
      20'h0dca8: out <= 12'h603;
      20'h0dca9: out <= 12'h603;
      20'h0dcaa: out <= 12'h603;
      20'h0dcab: out <= 12'h603;
      20'h0dcac: out <= 12'h603;
      20'h0dcad: out <= 12'h603;
      20'h0dcae: out <= 12'h603;
      20'h0dcaf: out <= 12'h603;
      20'h0dcb0: out <= 12'hee9;
      20'h0dcb1: out <= 12'hf87;
      20'h0dcb2: out <= 12'hf87;
      20'h0dcb3: out <= 12'hf87;
      20'h0dcb4: out <= 12'hf87;
      20'h0dcb5: out <= 12'hf87;
      20'h0dcb6: out <= 12'hf87;
      20'h0dcb7: out <= 12'hb27;
      20'h0dcb8: out <= 12'h000;
      20'h0dcb9: out <= 12'h000;
      20'h0dcba: out <= 12'h000;
      20'h0dcbb: out <= 12'h000;
      20'h0dcbc: out <= 12'h000;
      20'h0dcbd: out <= 12'h000;
      20'h0dcbe: out <= 12'h000;
      20'h0dcbf: out <= 12'h000;
      20'h0dcc0: out <= 12'h000;
      20'h0dcc1: out <= 12'h000;
      20'h0dcc2: out <= 12'h000;
      20'h0dcc3: out <= 12'h000;
      20'h0dcc4: out <= 12'h000;
      20'h0dcc5: out <= 12'h000;
      20'h0dcc6: out <= 12'h666;
      20'h0dcc7: out <= 12'hbbb;
      20'h0dcc8: out <= 12'hfff;
      20'h0dcc9: out <= 12'hbbb;
      20'h0dcca: out <= 12'h666;
      20'h0dccb: out <= 12'h000;
      20'h0dccc: out <= 12'h000;
      20'h0dccd: out <= 12'h000;
      20'h0dcce: out <= 12'h000;
      20'h0dccf: out <= 12'h000;
      20'h0dcd0: out <= 12'h000;
      20'h0dcd1: out <= 12'h000;
      20'h0dcd2: out <= 12'h000;
      20'h0dcd3: out <= 12'h000;
      20'h0dcd4: out <= 12'h000;
      20'h0dcd5: out <= 12'h000;
      20'h0dcd6: out <= 12'h000;
      20'h0dcd7: out <= 12'h000;
      20'h0dcd8: out <= 12'h000;
      20'h0dcd9: out <= 12'h000;
      20'h0dcda: out <= 12'h000;
      20'h0dcdb: out <= 12'h000;
      20'h0dcdc: out <= 12'h000;
      20'h0dcdd: out <= 12'h000;
      20'h0dcde: out <= 12'h000;
      20'h0dcdf: out <= 12'h000;
      20'h0dce0: out <= 12'h000;
      20'h0dce1: out <= 12'h000;
      20'h0dce2: out <= 12'h000;
      20'h0dce3: out <= 12'h000;
      20'h0dce4: out <= 12'h000;
      20'h0dce5: out <= 12'h000;
      20'h0dce6: out <= 12'h000;
      20'h0dce7: out <= 12'h000;
      20'h0dce8: out <= 12'h000;
      20'h0dce9: out <= 12'h000;
      20'h0dcea: out <= 12'h000;
      20'h0dceb: out <= 12'h000;
      20'h0dcec: out <= 12'h000;
      20'h0dced: out <= 12'h000;
      20'h0dcee: out <= 12'h000;
      20'h0dcef: out <= 12'h000;
      20'h0dcf0: out <= 12'h000;
      20'h0dcf1: out <= 12'hc7f;
      20'h0dcf2: out <= 12'hfff;
      20'h0dcf3: out <= 12'hfff;
      20'h0dcf4: out <= 12'h72f;
      20'h0dcf5: out <= 12'hc7f;
      20'h0dcf6: out <= 12'hfff;
      20'h0dcf7: out <= 12'hfff;
      20'h0dcf8: out <= 12'hfff;
      20'h0dcf9: out <= 12'hfff;
      20'h0dcfa: out <= 12'hc7f;
      20'h0dcfb: out <= 12'h72f;
      20'h0dcfc: out <= 12'hfff;
      20'h0dcfd: out <= 12'hfff;
      20'h0dcfe: out <= 12'hc7f;
      20'h0dcff: out <= 12'h000;
      20'h0dd00: out <= 12'h000;
      20'h0dd01: out <= 12'hbbb;
      20'h0dd02: out <= 12'hfff;
      20'h0dd03: out <= 12'h666;
      20'h0dd04: out <= 12'hbbb;
      20'h0dd05: out <= 12'hbbb;
      20'h0dd06: out <= 12'hbbb;
      20'h0dd07: out <= 12'h666;
      20'h0dd08: out <= 12'h666;
      20'h0dd09: out <= 12'h666;
      20'h0dd0a: out <= 12'h666;
      20'h0dd0b: out <= 12'h666;
      20'h0dd0c: out <= 12'h666;
      20'h0dd0d: out <= 12'hfff;
      20'h0dd0e: out <= 12'hbbb;
      20'h0dd0f: out <= 12'h000;
      20'h0dd10: out <= 12'h000;
      20'h0dd11: out <= 12'hbb0;
      20'h0dd12: out <= 12'hee9;
      20'h0dd13: out <= 12'hbb0;
      20'h0dd14: out <= 12'hbb0;
      20'h0dd15: out <= 12'h660;
      20'h0dd16: out <= 12'hbb0;
      20'h0dd17: out <= 12'hee9;
      20'h0dd18: out <= 12'hee9;
      20'h0dd19: out <= 12'hbb0;
      20'h0dd1a: out <= 12'h660;
      20'h0dd1b: out <= 12'hbb0;
      20'h0dd1c: out <= 12'hbb0;
      20'h0dd1d: out <= 12'hee9;
      20'h0dd1e: out <= 12'hbb0;
      20'h0dd1f: out <= 12'h000;
      20'h0dd20: out <= 12'h000;
      20'h0dd21: out <= 12'h6af;
      20'h0dd22: out <= 12'hfff;
      20'h0dd23: out <= 12'hfff;
      20'h0dd24: out <= 12'h6af;
      20'h0dd25: out <= 12'h16d;
      20'h0dd26: out <= 12'h16d;
      20'h0dd27: out <= 12'h16d;
      20'h0dd28: out <= 12'h16d;
      20'h0dd29: out <= 12'h16d;
      20'h0dd2a: out <= 12'h16d;
      20'h0dd2b: out <= 12'hfff;
      20'h0dd2c: out <= 12'hfff;
      20'h0dd2d: out <= 12'hfff;
      20'h0dd2e: out <= 12'h6af;
      20'h0dd2f: out <= 12'h000;
      20'h0dd30: out <= 12'h000;
      20'h0dd31: out <= 12'hc7f;
      20'h0dd32: out <= 12'hfff;
      20'h0dd33: out <= 12'h72f;
      20'h0dd34: out <= 12'hfff;
      20'h0dd35: out <= 12'hfff;
      20'h0dd36: out <= 12'hfff;
      20'h0dd37: out <= 12'h72f;
      20'h0dd38: out <= 12'h72f;
      20'h0dd39: out <= 12'hfff;
      20'h0dd3a: out <= 12'hfff;
      20'h0dd3b: out <= 12'hfff;
      20'h0dd3c: out <= 12'h72f;
      20'h0dd3d: out <= 12'hfff;
      20'h0dd3e: out <= 12'hc7f;
      20'h0dd3f: out <= 12'h000;
      20'h0dd40: out <= 12'h000;
      20'h0dd41: out <= 12'hbbb;
      20'h0dd42: out <= 12'hfff;
      20'h0dd43: out <= 12'hfff;
      20'h0dd44: out <= 12'hfff;
      20'h0dd45: out <= 12'h666;
      20'h0dd46: out <= 12'hbbb;
      20'h0dd47: out <= 12'hfff;
      20'h0dd48: out <= 12'hfff;
      20'h0dd49: out <= 12'hfff;
      20'h0dd4a: out <= 12'hfff;
      20'h0dd4b: out <= 12'hfff;
      20'h0dd4c: out <= 12'hfff;
      20'h0dd4d: out <= 12'hfff;
      20'h0dd4e: out <= 12'hbbb;
      20'h0dd4f: out <= 12'h000;
      20'h0dd50: out <= 12'h000;
      20'h0dd51: out <= 12'h6af;
      20'h0dd52: out <= 12'hfff;
      20'h0dd53: out <= 12'hfff;
      20'h0dd54: out <= 12'hfff;
      20'h0dd55: out <= 12'h6af;
      20'h0dd56: out <= 12'h6af;
      20'h0dd57: out <= 12'h16d;
      20'h0dd58: out <= 12'h6af;
      20'h0dd59: out <= 12'h16d;
      20'h0dd5a: out <= 12'h16d;
      20'h0dd5b: out <= 12'hfff;
      20'h0dd5c: out <= 12'hfff;
      20'h0dd5d: out <= 12'hfff;
      20'h0dd5e: out <= 12'h6af;
      20'h0dd5f: out <= 12'h000;
      20'h0dd60: out <= 12'h000;
      20'h0dd61: out <= 12'hbb0;
      20'h0dd62: out <= 12'hee9;
      20'h0dd63: out <= 12'hee9;
      20'h0dd64: out <= 12'hee9;
      20'h0dd65: out <= 12'h660;
      20'h0dd66: out <= 12'hbb0;
      20'h0dd67: out <= 12'hbb0;
      20'h0dd68: out <= 12'hbb0;
      20'h0dd69: out <= 12'hbb0;
      20'h0dd6a: out <= 12'h660;
      20'h0dd6b: out <= 12'hee9;
      20'h0dd6c: out <= 12'hee9;
      20'h0dd6d: out <= 12'hee9;
      20'h0dd6e: out <= 12'hbb0;
      20'h0dd6f: out <= 12'h000;
      20'h0dd70: out <= 12'h603;
      20'h0dd71: out <= 12'h603;
      20'h0dd72: out <= 12'h603;
      20'h0dd73: out <= 12'h603;
      20'h0dd74: out <= 12'h603;
      20'h0dd75: out <= 12'h603;
      20'h0dd76: out <= 12'h603;
      20'h0dd77: out <= 12'h603;
      20'h0dd78: out <= 12'h603;
      20'h0dd79: out <= 12'h603;
      20'h0dd7a: out <= 12'h603;
      20'h0dd7b: out <= 12'h603;
      20'h0dd7c: out <= 12'h603;
      20'h0dd7d: out <= 12'h603;
      20'h0dd7e: out <= 12'h603;
      20'h0dd7f: out <= 12'h603;
      20'h0dd80: out <= 12'h603;
      20'h0dd81: out <= 12'h603;
      20'h0dd82: out <= 12'h603;
      20'h0dd83: out <= 12'h603;
      20'h0dd84: out <= 12'h603;
      20'h0dd85: out <= 12'h603;
      20'h0dd86: out <= 12'h603;
      20'h0dd87: out <= 12'h603;
      20'h0dd88: out <= 12'h603;
      20'h0dd89: out <= 12'h603;
      20'h0dd8a: out <= 12'h603;
      20'h0dd8b: out <= 12'h603;
      20'h0dd8c: out <= 12'h603;
      20'h0dd8d: out <= 12'h603;
      20'h0dd8e: out <= 12'h603;
      20'h0dd8f: out <= 12'h603;
      20'h0dd90: out <= 12'h603;
      20'h0dd91: out <= 12'h603;
      20'h0dd92: out <= 12'h603;
      20'h0dd93: out <= 12'h603;
      20'h0dd94: out <= 12'h603;
      20'h0dd95: out <= 12'h603;
      20'h0dd96: out <= 12'h603;
      20'h0dd97: out <= 12'h603;
      20'h0dd98: out <= 12'h603;
      20'h0dd99: out <= 12'h603;
      20'h0dd9a: out <= 12'h603;
      20'h0dd9b: out <= 12'h603;
      20'h0dd9c: out <= 12'h603;
      20'h0dd9d: out <= 12'h603;
      20'h0dd9e: out <= 12'h603;
      20'h0dd9f: out <= 12'h603;
      20'h0dda0: out <= 12'h603;
      20'h0dda1: out <= 12'h603;
      20'h0dda2: out <= 12'h603;
      20'h0dda3: out <= 12'h603;
      20'h0dda4: out <= 12'h603;
      20'h0dda5: out <= 12'h603;
      20'h0dda6: out <= 12'h603;
      20'h0dda7: out <= 12'h603;
      20'h0dda8: out <= 12'h603;
      20'h0dda9: out <= 12'h603;
      20'h0ddaa: out <= 12'h603;
      20'h0ddab: out <= 12'h603;
      20'h0ddac: out <= 12'h603;
      20'h0ddad: out <= 12'h603;
      20'h0ddae: out <= 12'h603;
      20'h0ddaf: out <= 12'h603;
      20'h0ddb0: out <= 12'h603;
      20'h0ddb1: out <= 12'h603;
      20'h0ddb2: out <= 12'h603;
      20'h0ddb3: out <= 12'h603;
      20'h0ddb4: out <= 12'h603;
      20'h0ddb5: out <= 12'h603;
      20'h0ddb6: out <= 12'h603;
      20'h0ddb7: out <= 12'h603;
      20'h0ddb8: out <= 12'h603;
      20'h0ddb9: out <= 12'h603;
      20'h0ddba: out <= 12'h603;
      20'h0ddbb: out <= 12'h603;
      20'h0ddbc: out <= 12'h603;
      20'h0ddbd: out <= 12'h603;
      20'h0ddbe: out <= 12'h603;
      20'h0ddbf: out <= 12'h603;
      20'h0ddc0: out <= 12'h603;
      20'h0ddc1: out <= 12'h603;
      20'h0ddc2: out <= 12'h603;
      20'h0ddc3: out <= 12'h603;
      20'h0ddc4: out <= 12'h603;
      20'h0ddc5: out <= 12'h603;
      20'h0ddc6: out <= 12'h603;
      20'h0ddc7: out <= 12'h603;
      20'h0ddc8: out <= 12'hee9;
      20'h0ddc9: out <= 12'hf87;
      20'h0ddca: out <= 12'hee9;
      20'h0ddcb: out <= 12'hee9;
      20'h0ddcc: out <= 12'hee9;
      20'h0ddcd: out <= 12'hb27;
      20'h0ddce: out <= 12'hf87;
      20'h0ddcf: out <= 12'hb27;
      20'h0ddd0: out <= 12'h000;
      20'h0ddd1: out <= 12'h000;
      20'h0ddd2: out <= 12'h000;
      20'h0ddd3: out <= 12'h000;
      20'h0ddd4: out <= 12'h000;
      20'h0ddd5: out <= 12'h000;
      20'h0ddd6: out <= 12'h000;
      20'h0ddd7: out <= 12'h000;
      20'h0ddd8: out <= 12'h000;
      20'h0ddd9: out <= 12'h000;
      20'h0ddda: out <= 12'h000;
      20'h0dddb: out <= 12'h000;
      20'h0dddc: out <= 12'h000;
      20'h0dddd: out <= 12'h000;
      20'h0ddde: out <= 12'h666;
      20'h0dddf: out <= 12'hbbb;
      20'h0dde0: out <= 12'hfff;
      20'h0dde1: out <= 12'hbbb;
      20'h0dde2: out <= 12'h666;
      20'h0dde3: out <= 12'h000;
      20'h0dde4: out <= 12'h000;
      20'h0dde5: out <= 12'h000;
      20'h0dde6: out <= 12'h000;
      20'h0dde7: out <= 12'h000;
      20'h0dde8: out <= 12'h000;
      20'h0dde9: out <= 12'h000;
      20'h0ddea: out <= 12'h000;
      20'h0ddeb: out <= 12'h000;
      20'h0ddec: out <= 12'h000;
      20'h0dded: out <= 12'h000;
      20'h0ddee: out <= 12'h000;
      20'h0ddef: out <= 12'h000;
      20'h0ddf0: out <= 12'h000;
      20'h0ddf1: out <= 12'h000;
      20'h0ddf2: out <= 12'h000;
      20'h0ddf3: out <= 12'h000;
      20'h0ddf4: out <= 12'h000;
      20'h0ddf5: out <= 12'h000;
      20'h0ddf6: out <= 12'h000;
      20'h0ddf7: out <= 12'h000;
      20'h0ddf8: out <= 12'h000;
      20'h0ddf9: out <= 12'h000;
      20'h0ddfa: out <= 12'h000;
      20'h0ddfb: out <= 12'h000;
      20'h0ddfc: out <= 12'h000;
      20'h0ddfd: out <= 12'h000;
      20'h0ddfe: out <= 12'h000;
      20'h0ddff: out <= 12'h000;
      20'h0de00: out <= 12'h000;
      20'h0de01: out <= 12'h000;
      20'h0de02: out <= 12'h000;
      20'h0de03: out <= 12'h000;
      20'h0de04: out <= 12'h000;
      20'h0de05: out <= 12'h000;
      20'h0de06: out <= 12'h000;
      20'h0de07: out <= 12'h000;
      20'h0de08: out <= 12'h000;
      20'h0de09: out <= 12'h72f;
      20'h0de0a: out <= 12'hfff;
      20'h0de0b: out <= 12'hfff;
      20'h0de0c: out <= 12'hc7f;
      20'h0de0d: out <= 12'h72f;
      20'h0de0e: out <= 12'hc7f;
      20'h0de0f: out <= 12'hc7f;
      20'h0de10: out <= 12'hc7f;
      20'h0de11: out <= 12'hc7f;
      20'h0de12: out <= 12'h72f;
      20'h0de13: out <= 12'hc7f;
      20'h0de14: out <= 12'hfff;
      20'h0de15: out <= 12'hfff;
      20'h0de16: out <= 12'h72f;
      20'h0de17: out <= 12'h000;
      20'h0de18: out <= 12'h000;
      20'h0de19: out <= 12'h666;
      20'h0de1a: out <= 12'hfff;
      20'h0de1b: out <= 12'hfff;
      20'h0de1c: out <= 12'h666;
      20'h0de1d: out <= 12'hbbb;
      20'h0de1e: out <= 12'hbbb;
      20'h0de1f: out <= 12'h666;
      20'h0de20: out <= 12'h666;
      20'h0de21: out <= 12'h666;
      20'h0de22: out <= 12'h666;
      20'h0de23: out <= 12'h666;
      20'h0de24: out <= 12'hfff;
      20'h0de25: out <= 12'hfff;
      20'h0de26: out <= 12'h666;
      20'h0de27: out <= 12'h000;
      20'h0de28: out <= 12'h000;
      20'h0de29: out <= 12'h660;
      20'h0de2a: out <= 12'hee9;
      20'h0de2b: out <= 12'h660;
      20'h0de2c: out <= 12'h660;
      20'h0de2d: out <= 12'h660;
      20'h0de2e: out <= 12'h660;
      20'h0de2f: out <= 12'h660;
      20'h0de30: out <= 12'h660;
      20'h0de31: out <= 12'h660;
      20'h0de32: out <= 12'h660;
      20'h0de33: out <= 12'h660;
      20'h0de34: out <= 12'h660;
      20'h0de35: out <= 12'hee9;
      20'h0de36: out <= 12'h660;
      20'h0de37: out <= 12'h000;
      20'h0de38: out <= 12'h000;
      20'h0de39: out <= 12'h16d;
      20'h0de3a: out <= 12'hfff;
      20'h0de3b: out <= 12'hfff;
      20'h0de3c: out <= 12'h6af;
      20'h0de3d: out <= 12'h16d;
      20'h0de3e: out <= 12'h16d;
      20'h0de3f: out <= 12'hfff;
      20'h0de40: out <= 12'hfff;
      20'h0de41: out <= 12'hfff;
      20'h0de42: out <= 12'hfff;
      20'h0de43: out <= 12'hfff;
      20'h0de44: out <= 12'hfff;
      20'h0de45: out <= 12'hfff;
      20'h0de46: out <= 12'h16d;
      20'h0de47: out <= 12'h000;
      20'h0de48: out <= 12'h000;
      20'h0de49: out <= 12'h72f;
      20'h0de4a: out <= 12'hfff;
      20'h0de4b: out <= 12'hfff;
      20'h0de4c: out <= 12'hfff;
      20'h0de4d: out <= 12'hfff;
      20'h0de4e: out <= 12'hfff;
      20'h0de4f: out <= 12'hc7f;
      20'h0de50: out <= 12'hc7f;
      20'h0de51: out <= 12'hfff;
      20'h0de52: out <= 12'hfff;
      20'h0de53: out <= 12'hfff;
      20'h0de54: out <= 12'hfff;
      20'h0de55: out <= 12'hfff;
      20'h0de56: out <= 12'h72f;
      20'h0de57: out <= 12'h000;
      20'h0de58: out <= 12'h000;
      20'h0de59: out <= 12'h666;
      20'h0de5a: out <= 12'hfff;
      20'h0de5b: out <= 12'hfff;
      20'h0de5c: out <= 12'h666;
      20'h0de5d: out <= 12'hbbb;
      20'h0de5e: out <= 12'h666;
      20'h0de5f: out <= 12'hbbb;
      20'h0de60: out <= 12'hbbb;
      20'h0de61: out <= 12'h666;
      20'h0de62: out <= 12'h666;
      20'h0de63: out <= 12'hfff;
      20'h0de64: out <= 12'hfff;
      20'h0de65: out <= 12'hfff;
      20'h0de66: out <= 12'h666;
      20'h0de67: out <= 12'h000;
      20'h0de68: out <= 12'h000;
      20'h0de69: out <= 12'h16d;
      20'h0de6a: out <= 12'hfff;
      20'h0de6b: out <= 12'hfff;
      20'h0de6c: out <= 12'h16d;
      20'h0de6d: out <= 12'h6af;
      20'h0de6e: out <= 12'h6af;
      20'h0de6f: out <= 12'h16d;
      20'h0de70: out <= 12'h6af;
      20'h0de71: out <= 12'h16d;
      20'h0de72: out <= 12'h16d;
      20'h0de73: out <= 12'h16d;
      20'h0de74: out <= 12'hfff;
      20'h0de75: out <= 12'hfff;
      20'h0de76: out <= 12'h16d;
      20'h0de77: out <= 12'h000;
      20'h0de78: out <= 12'h000;
      20'h0de79: out <= 12'h660;
      20'h0de7a: out <= 12'hee9;
      20'h0de7b: out <= 12'hee9;
      20'h0de7c: out <= 12'hee9;
      20'h0de7d: out <= 12'hee9;
      20'h0de7e: out <= 12'h660;
      20'h0de7f: out <= 12'hbb0;
      20'h0de80: out <= 12'hbb0;
      20'h0de81: out <= 12'h660;
      20'h0de82: out <= 12'hee9;
      20'h0de83: out <= 12'hee9;
      20'h0de84: out <= 12'hee9;
      20'h0de85: out <= 12'hee9;
      20'h0de86: out <= 12'h660;
      20'h0de87: out <= 12'h000;
      20'h0de88: out <= 12'h603;
      20'h0de89: out <= 12'h603;
      20'h0de8a: out <= 12'h603;
      20'h0de8b: out <= 12'h603;
      20'h0de8c: out <= 12'h603;
      20'h0de8d: out <= 12'h603;
      20'h0de8e: out <= 12'h603;
      20'h0de8f: out <= 12'h603;
      20'h0de90: out <= 12'h603;
      20'h0de91: out <= 12'h603;
      20'h0de92: out <= 12'h603;
      20'h0de93: out <= 12'h603;
      20'h0de94: out <= 12'h603;
      20'h0de95: out <= 12'h603;
      20'h0de96: out <= 12'h603;
      20'h0de97: out <= 12'h603;
      20'h0de98: out <= 12'h603;
      20'h0de99: out <= 12'h603;
      20'h0de9a: out <= 12'h603;
      20'h0de9b: out <= 12'h603;
      20'h0de9c: out <= 12'h603;
      20'h0de9d: out <= 12'h603;
      20'h0de9e: out <= 12'h603;
      20'h0de9f: out <= 12'h603;
      20'h0dea0: out <= 12'h603;
      20'h0dea1: out <= 12'h603;
      20'h0dea2: out <= 12'h603;
      20'h0dea3: out <= 12'h603;
      20'h0dea4: out <= 12'h603;
      20'h0dea5: out <= 12'h603;
      20'h0dea6: out <= 12'h603;
      20'h0dea7: out <= 12'h603;
      20'h0dea8: out <= 12'h603;
      20'h0dea9: out <= 12'h603;
      20'h0deaa: out <= 12'h603;
      20'h0deab: out <= 12'h603;
      20'h0deac: out <= 12'h603;
      20'h0dead: out <= 12'h603;
      20'h0deae: out <= 12'h603;
      20'h0deaf: out <= 12'h603;
      20'h0deb0: out <= 12'h603;
      20'h0deb1: out <= 12'h603;
      20'h0deb2: out <= 12'h603;
      20'h0deb3: out <= 12'h603;
      20'h0deb4: out <= 12'h603;
      20'h0deb5: out <= 12'h603;
      20'h0deb6: out <= 12'h603;
      20'h0deb7: out <= 12'h603;
      20'h0deb8: out <= 12'h603;
      20'h0deb9: out <= 12'h603;
      20'h0deba: out <= 12'h603;
      20'h0debb: out <= 12'h603;
      20'h0debc: out <= 12'h603;
      20'h0debd: out <= 12'h603;
      20'h0debe: out <= 12'h603;
      20'h0debf: out <= 12'h603;
      20'h0dec0: out <= 12'h603;
      20'h0dec1: out <= 12'h603;
      20'h0dec2: out <= 12'h603;
      20'h0dec3: out <= 12'h603;
      20'h0dec4: out <= 12'h603;
      20'h0dec5: out <= 12'h603;
      20'h0dec6: out <= 12'h603;
      20'h0dec7: out <= 12'h603;
      20'h0dec8: out <= 12'h603;
      20'h0dec9: out <= 12'h603;
      20'h0deca: out <= 12'h603;
      20'h0decb: out <= 12'h603;
      20'h0decc: out <= 12'h603;
      20'h0decd: out <= 12'h603;
      20'h0dece: out <= 12'h603;
      20'h0decf: out <= 12'h603;
      20'h0ded0: out <= 12'h603;
      20'h0ded1: out <= 12'h603;
      20'h0ded2: out <= 12'h603;
      20'h0ded3: out <= 12'h603;
      20'h0ded4: out <= 12'h603;
      20'h0ded5: out <= 12'h603;
      20'h0ded6: out <= 12'h603;
      20'h0ded7: out <= 12'h603;
      20'h0ded8: out <= 12'h603;
      20'h0ded9: out <= 12'h603;
      20'h0deda: out <= 12'h603;
      20'h0dedb: out <= 12'h603;
      20'h0dedc: out <= 12'h603;
      20'h0dedd: out <= 12'h603;
      20'h0dede: out <= 12'h603;
      20'h0dedf: out <= 12'h603;
      20'h0dee0: out <= 12'hee9;
      20'h0dee1: out <= 12'hf87;
      20'h0dee2: out <= 12'hee9;
      20'h0dee3: out <= 12'hf87;
      20'h0dee4: out <= 12'hf87;
      20'h0dee5: out <= 12'hb27;
      20'h0dee6: out <= 12'hf87;
      20'h0dee7: out <= 12'hb27;
      20'h0dee8: out <= 12'h000;
      20'h0dee9: out <= 12'h000;
      20'h0deea: out <= 12'h000;
      20'h0deeb: out <= 12'h000;
      20'h0deec: out <= 12'h000;
      20'h0deed: out <= 12'h000;
      20'h0deee: out <= 12'h000;
      20'h0deef: out <= 12'h000;
      20'h0def0: out <= 12'h000;
      20'h0def1: out <= 12'h000;
      20'h0def2: out <= 12'h000;
      20'h0def3: out <= 12'hbbb;
      20'h0def4: out <= 12'h000;
      20'h0def5: out <= 12'h666;
      20'h0def6: out <= 12'h666;
      20'h0def7: out <= 12'hbbb;
      20'h0def8: out <= 12'hfff;
      20'h0def9: out <= 12'hbbb;
      20'h0defa: out <= 12'h666;
      20'h0defb: out <= 12'h666;
      20'h0defc: out <= 12'h000;
      20'h0defd: out <= 12'hbbb;
      20'h0defe: out <= 12'h000;
      20'h0deff: out <= 12'h000;
      20'h0df00: out <= 12'h000;
      20'h0df01: out <= 12'h000;
      20'h0df02: out <= 12'h000;
      20'h0df03: out <= 12'h000;
      20'h0df04: out <= 12'h000;
      20'h0df05: out <= 12'h000;
      20'h0df06: out <= 12'h000;
      20'h0df07: out <= 12'h000;
      20'h0df08: out <= 12'h000;
      20'h0df09: out <= 12'h000;
      20'h0df0a: out <= 12'h000;
      20'h0df0b: out <= 12'h000;
      20'h0df0c: out <= 12'h000;
      20'h0df0d: out <= 12'h000;
      20'h0df0e: out <= 12'h000;
      20'h0df0f: out <= 12'h000;
      20'h0df10: out <= 12'h000;
      20'h0df11: out <= 12'h000;
      20'h0df12: out <= 12'h000;
      20'h0df13: out <= 12'h000;
      20'h0df14: out <= 12'h000;
      20'h0df15: out <= 12'h000;
      20'h0df16: out <= 12'h000;
      20'h0df17: out <= 12'h000;
      20'h0df18: out <= 12'h000;
      20'h0df19: out <= 12'h000;
      20'h0df1a: out <= 12'h000;
      20'h0df1b: out <= 12'h000;
      20'h0df1c: out <= 12'h000;
      20'h0df1d: out <= 12'h000;
      20'h0df1e: out <= 12'h000;
      20'h0df1f: out <= 12'h000;
      20'h0df20: out <= 12'h000;
      20'h0df21: out <= 12'h72f;
      20'h0df22: out <= 12'hfff;
      20'h0df23: out <= 12'hfff;
      20'h0df24: out <= 12'hfff;
      20'h0df25: out <= 12'hfff;
      20'h0df26: out <= 12'h72f;
      20'h0df27: out <= 12'h72f;
      20'h0df28: out <= 12'h72f;
      20'h0df29: out <= 12'h72f;
      20'h0df2a: out <= 12'hfff;
      20'h0df2b: out <= 12'hfff;
      20'h0df2c: out <= 12'hfff;
      20'h0df2d: out <= 12'hfff;
      20'h0df2e: out <= 12'h72f;
      20'h0df2f: out <= 12'h000;
      20'h0df30: out <= 12'h000;
      20'h0df31: out <= 12'h666;
      20'h0df32: out <= 12'hfff;
      20'h0df33: out <= 12'hfff;
      20'h0df34: out <= 12'hfff;
      20'h0df35: out <= 12'h666;
      20'h0df36: out <= 12'h666;
      20'h0df37: out <= 12'h666;
      20'h0df38: out <= 12'h666;
      20'h0df39: out <= 12'h666;
      20'h0df3a: out <= 12'h666;
      20'h0df3b: out <= 12'hfff;
      20'h0df3c: out <= 12'hfff;
      20'h0df3d: out <= 12'hfff;
      20'h0df3e: out <= 12'h666;
      20'h0df3f: out <= 12'h000;
      20'h0df40: out <= 12'h000;
      20'h0df41: out <= 12'h660;
      20'h0df42: out <= 12'hee9;
      20'h0df43: out <= 12'hbb0;
      20'h0df44: out <= 12'hbb0;
      20'h0df45: out <= 12'hee9;
      20'h0df46: out <= 12'hee9;
      20'h0df47: out <= 12'hee9;
      20'h0df48: out <= 12'hee9;
      20'h0df49: out <= 12'hee9;
      20'h0df4a: out <= 12'hee9;
      20'h0df4b: out <= 12'hbb0;
      20'h0df4c: out <= 12'hbb0;
      20'h0df4d: out <= 12'hee9;
      20'h0df4e: out <= 12'h660;
      20'h0df4f: out <= 12'h000;
      20'h0df50: out <= 12'h000;
      20'h0df51: out <= 12'h16d;
      20'h0df52: out <= 12'hfff;
      20'h0df53: out <= 12'hfff;
      20'h0df54: out <= 12'h6af;
      20'h0df55: out <= 12'h16d;
      20'h0df56: out <= 12'h16d;
      20'h0df57: out <= 12'hfff;
      20'h0df58: out <= 12'hfff;
      20'h0df59: out <= 12'hfff;
      20'h0df5a: out <= 12'hfff;
      20'h0df5b: out <= 12'hfff;
      20'h0df5c: out <= 12'hfff;
      20'h0df5d: out <= 12'hfff;
      20'h0df5e: out <= 12'h16d;
      20'h0df5f: out <= 12'h000;
      20'h0df60: out <= 12'h000;
      20'h0df61: out <= 12'h72f;
      20'h0df62: out <= 12'hfff;
      20'h0df63: out <= 12'hfff;
      20'h0df64: out <= 12'hfff;
      20'h0df65: out <= 12'hfff;
      20'h0df66: out <= 12'h72f;
      20'h0df67: out <= 12'hc7f;
      20'h0df68: out <= 12'hc7f;
      20'h0df69: out <= 12'h72f;
      20'h0df6a: out <= 12'hfff;
      20'h0df6b: out <= 12'hfff;
      20'h0df6c: out <= 12'hfff;
      20'h0df6d: out <= 12'hfff;
      20'h0df6e: out <= 12'h72f;
      20'h0df6f: out <= 12'h000;
      20'h0df70: out <= 12'h000;
      20'h0df71: out <= 12'h666;
      20'h0df72: out <= 12'hfff;
      20'h0df73: out <= 12'hfff;
      20'h0df74: out <= 12'h666;
      20'h0df75: out <= 12'hbbb;
      20'h0df76: out <= 12'h666;
      20'h0df77: out <= 12'hbbb;
      20'h0df78: out <= 12'hbbb;
      20'h0df79: out <= 12'h666;
      20'h0df7a: out <= 12'h666;
      20'h0df7b: out <= 12'hfff;
      20'h0df7c: out <= 12'hfff;
      20'h0df7d: out <= 12'hfff;
      20'h0df7e: out <= 12'h666;
      20'h0df7f: out <= 12'h000;
      20'h0df80: out <= 12'h000;
      20'h0df81: out <= 12'h16d;
      20'h0df82: out <= 12'hfff;
      20'h0df83: out <= 12'hfff;
      20'h0df84: out <= 12'h16d;
      20'h0df85: out <= 12'h6af;
      20'h0df86: out <= 12'h6af;
      20'h0df87: out <= 12'h16d;
      20'h0df88: out <= 12'h6af;
      20'h0df89: out <= 12'h16d;
      20'h0df8a: out <= 12'h16d;
      20'h0df8b: out <= 12'h16d;
      20'h0df8c: out <= 12'hfff;
      20'h0df8d: out <= 12'hfff;
      20'h0df8e: out <= 12'h16d;
      20'h0df8f: out <= 12'h000;
      20'h0df90: out <= 12'h000;
      20'h0df91: out <= 12'h660;
      20'h0df92: out <= 12'hee9;
      20'h0df93: out <= 12'hee9;
      20'h0df94: out <= 12'hee9;
      20'h0df95: out <= 12'hee9;
      20'h0df96: out <= 12'hee9;
      20'h0df97: out <= 12'h660;
      20'h0df98: out <= 12'h660;
      20'h0df99: out <= 12'hee9;
      20'h0df9a: out <= 12'hee9;
      20'h0df9b: out <= 12'hee9;
      20'h0df9c: out <= 12'hee9;
      20'h0df9d: out <= 12'hee9;
      20'h0df9e: out <= 12'h660;
      20'h0df9f: out <= 12'h000;
      20'h0dfa0: out <= 12'h603;
      20'h0dfa1: out <= 12'h603;
      20'h0dfa2: out <= 12'h603;
      20'h0dfa3: out <= 12'h603;
      20'h0dfa4: out <= 12'h603;
      20'h0dfa5: out <= 12'h603;
      20'h0dfa6: out <= 12'h603;
      20'h0dfa7: out <= 12'h603;
      20'h0dfa8: out <= 12'h603;
      20'h0dfa9: out <= 12'h603;
      20'h0dfaa: out <= 12'h603;
      20'h0dfab: out <= 12'h603;
      20'h0dfac: out <= 12'h603;
      20'h0dfad: out <= 12'h603;
      20'h0dfae: out <= 12'h603;
      20'h0dfaf: out <= 12'h603;
      20'h0dfb0: out <= 12'h603;
      20'h0dfb1: out <= 12'h603;
      20'h0dfb2: out <= 12'h603;
      20'h0dfb3: out <= 12'h603;
      20'h0dfb4: out <= 12'h603;
      20'h0dfb5: out <= 12'h603;
      20'h0dfb6: out <= 12'h603;
      20'h0dfb7: out <= 12'h603;
      20'h0dfb8: out <= 12'h603;
      20'h0dfb9: out <= 12'h603;
      20'h0dfba: out <= 12'h603;
      20'h0dfbb: out <= 12'h603;
      20'h0dfbc: out <= 12'h603;
      20'h0dfbd: out <= 12'h603;
      20'h0dfbe: out <= 12'h603;
      20'h0dfbf: out <= 12'h603;
      20'h0dfc0: out <= 12'h603;
      20'h0dfc1: out <= 12'h603;
      20'h0dfc2: out <= 12'h603;
      20'h0dfc3: out <= 12'h603;
      20'h0dfc4: out <= 12'h603;
      20'h0dfc5: out <= 12'h603;
      20'h0dfc6: out <= 12'h603;
      20'h0dfc7: out <= 12'h603;
      20'h0dfc8: out <= 12'h603;
      20'h0dfc9: out <= 12'h603;
      20'h0dfca: out <= 12'h603;
      20'h0dfcb: out <= 12'h603;
      20'h0dfcc: out <= 12'h603;
      20'h0dfcd: out <= 12'h603;
      20'h0dfce: out <= 12'h603;
      20'h0dfcf: out <= 12'h603;
      20'h0dfd0: out <= 12'h603;
      20'h0dfd1: out <= 12'h603;
      20'h0dfd2: out <= 12'h603;
      20'h0dfd3: out <= 12'h603;
      20'h0dfd4: out <= 12'h603;
      20'h0dfd5: out <= 12'h603;
      20'h0dfd6: out <= 12'h603;
      20'h0dfd7: out <= 12'h603;
      20'h0dfd8: out <= 12'h603;
      20'h0dfd9: out <= 12'h603;
      20'h0dfda: out <= 12'h603;
      20'h0dfdb: out <= 12'h603;
      20'h0dfdc: out <= 12'h603;
      20'h0dfdd: out <= 12'h603;
      20'h0dfde: out <= 12'h603;
      20'h0dfdf: out <= 12'h603;
      20'h0dfe0: out <= 12'h603;
      20'h0dfe1: out <= 12'h603;
      20'h0dfe2: out <= 12'h603;
      20'h0dfe3: out <= 12'h603;
      20'h0dfe4: out <= 12'h603;
      20'h0dfe5: out <= 12'h603;
      20'h0dfe6: out <= 12'h603;
      20'h0dfe7: out <= 12'h603;
      20'h0dfe8: out <= 12'h603;
      20'h0dfe9: out <= 12'h603;
      20'h0dfea: out <= 12'h603;
      20'h0dfeb: out <= 12'h603;
      20'h0dfec: out <= 12'h603;
      20'h0dfed: out <= 12'h603;
      20'h0dfee: out <= 12'h603;
      20'h0dfef: out <= 12'h603;
      20'h0dff0: out <= 12'h603;
      20'h0dff1: out <= 12'h603;
      20'h0dff2: out <= 12'h603;
      20'h0dff3: out <= 12'h603;
      20'h0dff4: out <= 12'h603;
      20'h0dff5: out <= 12'h603;
      20'h0dff6: out <= 12'h603;
      20'h0dff7: out <= 12'h603;
      20'h0dff8: out <= 12'hee9;
      20'h0dff9: out <= 12'hf87;
      20'h0dffa: out <= 12'hee9;
      20'h0dffb: out <= 12'hf87;
      20'h0dffc: out <= 12'hf87;
      20'h0dffd: out <= 12'hb27;
      20'h0dffe: out <= 12'hf87;
      20'h0dfff: out <= 12'hb27;
      20'h0e000: out <= 12'h000;
      20'h0e001: out <= 12'h000;
      20'h0e002: out <= 12'h000;
      20'h0e003: out <= 12'h000;
      20'h0e004: out <= 12'h000;
      20'h0e005: out <= 12'h000;
      20'h0e006: out <= 12'h000;
      20'h0e007: out <= 12'h000;
      20'h0e008: out <= 12'h000;
      20'h0e009: out <= 12'h000;
      20'h0e00a: out <= 12'h666;
      20'h0e00b: out <= 12'hbbb;
      20'h0e00c: out <= 12'h666;
      20'h0e00d: out <= 12'hfff;
      20'h0e00e: out <= 12'h666;
      20'h0e00f: out <= 12'hbbb;
      20'h0e010: out <= 12'hfff;
      20'h0e011: out <= 12'hbbb;
      20'h0e012: out <= 12'h666;
      20'h0e013: out <= 12'h666;
      20'h0e014: out <= 12'h666;
      20'h0e015: out <= 12'hbbb;
      20'h0e016: out <= 12'h666;
      20'h0e017: out <= 12'h000;
      20'h0e018: out <= 12'h000;
      20'h0e019: out <= 12'h000;
      20'h0e01a: out <= 12'h000;
      20'h0e01b: out <= 12'h000;
      20'h0e01c: out <= 12'h000;
      20'h0e01d: out <= 12'h000;
      20'h0e01e: out <= 12'h000;
      20'h0e01f: out <= 12'h000;
      20'h0e020: out <= 12'h000;
      20'h0e021: out <= 12'h000;
      20'h0e022: out <= 12'h000;
      20'h0e023: out <= 12'h000;
      20'h0e024: out <= 12'h000;
      20'h0e025: out <= 12'h000;
      20'h0e026: out <= 12'h000;
      20'h0e027: out <= 12'h000;
      20'h0e028: out <= 12'h000;
      20'h0e029: out <= 12'h000;
      20'h0e02a: out <= 12'h000;
      20'h0e02b: out <= 12'h000;
      20'h0e02c: out <= 12'h000;
      20'h0e02d: out <= 12'h000;
      20'h0e02e: out <= 12'h000;
      20'h0e02f: out <= 12'h000;
      20'h0e030: out <= 12'h000;
      20'h0e031: out <= 12'h000;
      20'h0e032: out <= 12'h000;
      20'h0e033: out <= 12'h000;
      20'h0e034: out <= 12'h000;
      20'h0e035: out <= 12'h000;
      20'h0e036: out <= 12'h000;
      20'h0e037: out <= 12'h000;
      20'h0e038: out <= 12'h000;
      20'h0e039: out <= 12'h72f;
      20'h0e03a: out <= 12'h72f;
      20'h0e03b: out <= 12'hfff;
      20'h0e03c: out <= 12'hfff;
      20'h0e03d: out <= 12'hfff;
      20'h0e03e: out <= 12'hfff;
      20'h0e03f: out <= 12'hfff;
      20'h0e040: out <= 12'hfff;
      20'h0e041: out <= 12'hfff;
      20'h0e042: out <= 12'hfff;
      20'h0e043: out <= 12'hfff;
      20'h0e044: out <= 12'hfff;
      20'h0e045: out <= 12'h72f;
      20'h0e046: out <= 12'h72f;
      20'h0e047: out <= 12'h000;
      20'h0e048: out <= 12'h000;
      20'h0e049: out <= 12'h666;
      20'h0e04a: out <= 12'h666;
      20'h0e04b: out <= 12'hfff;
      20'h0e04c: out <= 12'hfff;
      20'h0e04d: out <= 12'hfff;
      20'h0e04e: out <= 12'hfff;
      20'h0e04f: out <= 12'hfff;
      20'h0e050: out <= 12'hfff;
      20'h0e051: out <= 12'hfff;
      20'h0e052: out <= 12'hfff;
      20'h0e053: out <= 12'hfff;
      20'h0e054: out <= 12'hfff;
      20'h0e055: out <= 12'h666;
      20'h0e056: out <= 12'h666;
      20'h0e057: out <= 12'h000;
      20'h0e058: out <= 12'h000;
      20'h0e059: out <= 12'h660;
      20'h0e05a: out <= 12'h660;
      20'h0e05b: out <= 12'hee9;
      20'h0e05c: out <= 12'hee9;
      20'h0e05d: out <= 12'hee9;
      20'h0e05e: out <= 12'hee9;
      20'h0e05f: out <= 12'hee9;
      20'h0e060: out <= 12'hee9;
      20'h0e061: out <= 12'hee9;
      20'h0e062: out <= 12'hee9;
      20'h0e063: out <= 12'hee9;
      20'h0e064: out <= 12'hee9;
      20'h0e065: out <= 12'h660;
      20'h0e066: out <= 12'h660;
      20'h0e067: out <= 12'h000;
      20'h0e068: out <= 12'h000;
      20'h0e069: out <= 12'h16d;
      20'h0e06a: out <= 12'h16d;
      20'h0e06b: out <= 12'hfff;
      20'h0e06c: out <= 12'hfff;
      20'h0e06d: out <= 12'hfff;
      20'h0e06e: out <= 12'hfff;
      20'h0e06f: out <= 12'hfff;
      20'h0e070: out <= 12'hfff;
      20'h0e071: out <= 12'hfff;
      20'h0e072: out <= 12'hfff;
      20'h0e073: out <= 12'hfff;
      20'h0e074: out <= 12'hfff;
      20'h0e075: out <= 12'h16d;
      20'h0e076: out <= 12'h16d;
      20'h0e077: out <= 12'h000;
      20'h0e078: out <= 12'h000;
      20'h0e079: out <= 12'h72f;
      20'h0e07a: out <= 12'h72f;
      20'h0e07b: out <= 12'hfff;
      20'h0e07c: out <= 12'hfff;
      20'h0e07d: out <= 12'hfff;
      20'h0e07e: out <= 12'hfff;
      20'h0e07f: out <= 12'hfff;
      20'h0e080: out <= 12'hfff;
      20'h0e081: out <= 12'hfff;
      20'h0e082: out <= 12'hfff;
      20'h0e083: out <= 12'hfff;
      20'h0e084: out <= 12'hfff;
      20'h0e085: out <= 12'h72f;
      20'h0e086: out <= 12'h72f;
      20'h0e087: out <= 12'h000;
      20'h0e088: out <= 12'h000;
      20'h0e089: out <= 12'h666;
      20'h0e08a: out <= 12'h666;
      20'h0e08b: out <= 12'hfff;
      20'h0e08c: out <= 12'hfff;
      20'h0e08d: out <= 12'hfff;
      20'h0e08e: out <= 12'hfff;
      20'h0e08f: out <= 12'hfff;
      20'h0e090: out <= 12'hfff;
      20'h0e091: out <= 12'hfff;
      20'h0e092: out <= 12'hfff;
      20'h0e093: out <= 12'hfff;
      20'h0e094: out <= 12'hfff;
      20'h0e095: out <= 12'h666;
      20'h0e096: out <= 12'h666;
      20'h0e097: out <= 12'h000;
      20'h0e098: out <= 12'h000;
      20'h0e099: out <= 12'h16d;
      20'h0e09a: out <= 12'h16d;
      20'h0e09b: out <= 12'hfff;
      20'h0e09c: out <= 12'hfff;
      20'h0e09d: out <= 12'hfff;
      20'h0e09e: out <= 12'hfff;
      20'h0e09f: out <= 12'hfff;
      20'h0e0a0: out <= 12'hfff;
      20'h0e0a1: out <= 12'hfff;
      20'h0e0a2: out <= 12'hfff;
      20'h0e0a3: out <= 12'hfff;
      20'h0e0a4: out <= 12'hfff;
      20'h0e0a5: out <= 12'h16d;
      20'h0e0a6: out <= 12'h16d;
      20'h0e0a7: out <= 12'h000;
      20'h0e0a8: out <= 12'h000;
      20'h0e0a9: out <= 12'h660;
      20'h0e0aa: out <= 12'h660;
      20'h0e0ab: out <= 12'hee9;
      20'h0e0ac: out <= 12'hee9;
      20'h0e0ad: out <= 12'hee9;
      20'h0e0ae: out <= 12'hee9;
      20'h0e0af: out <= 12'hee9;
      20'h0e0b0: out <= 12'hee9;
      20'h0e0b1: out <= 12'hee9;
      20'h0e0b2: out <= 12'hee9;
      20'h0e0b3: out <= 12'hee9;
      20'h0e0b4: out <= 12'hee9;
      20'h0e0b5: out <= 12'h660;
      20'h0e0b6: out <= 12'h660;
      20'h0e0b7: out <= 12'h000;
      20'h0e0b8: out <= 12'h603;
      20'h0e0b9: out <= 12'h603;
      20'h0e0ba: out <= 12'h603;
      20'h0e0bb: out <= 12'h603;
      20'h0e0bc: out <= 12'h603;
      20'h0e0bd: out <= 12'h603;
      20'h0e0be: out <= 12'h603;
      20'h0e0bf: out <= 12'h603;
      20'h0e0c0: out <= 12'h603;
      20'h0e0c1: out <= 12'h603;
      20'h0e0c2: out <= 12'h603;
      20'h0e0c3: out <= 12'h603;
      20'h0e0c4: out <= 12'h603;
      20'h0e0c5: out <= 12'h603;
      20'h0e0c6: out <= 12'h603;
      20'h0e0c7: out <= 12'h603;
      20'h0e0c8: out <= 12'h603;
      20'h0e0c9: out <= 12'h603;
      20'h0e0ca: out <= 12'h603;
      20'h0e0cb: out <= 12'h603;
      20'h0e0cc: out <= 12'h603;
      20'h0e0cd: out <= 12'h603;
      20'h0e0ce: out <= 12'h603;
      20'h0e0cf: out <= 12'h603;
      20'h0e0d0: out <= 12'h603;
      20'h0e0d1: out <= 12'h603;
      20'h0e0d2: out <= 12'h603;
      20'h0e0d3: out <= 12'h603;
      20'h0e0d4: out <= 12'h603;
      20'h0e0d5: out <= 12'h603;
      20'h0e0d6: out <= 12'h603;
      20'h0e0d7: out <= 12'h603;
      20'h0e0d8: out <= 12'h603;
      20'h0e0d9: out <= 12'h603;
      20'h0e0da: out <= 12'h603;
      20'h0e0db: out <= 12'h603;
      20'h0e0dc: out <= 12'h603;
      20'h0e0dd: out <= 12'h603;
      20'h0e0de: out <= 12'h603;
      20'h0e0df: out <= 12'h603;
      20'h0e0e0: out <= 12'h603;
      20'h0e0e1: out <= 12'h603;
      20'h0e0e2: out <= 12'h603;
      20'h0e0e3: out <= 12'h603;
      20'h0e0e4: out <= 12'h603;
      20'h0e0e5: out <= 12'h603;
      20'h0e0e6: out <= 12'h603;
      20'h0e0e7: out <= 12'h603;
      20'h0e0e8: out <= 12'h603;
      20'h0e0e9: out <= 12'h603;
      20'h0e0ea: out <= 12'h603;
      20'h0e0eb: out <= 12'h603;
      20'h0e0ec: out <= 12'h603;
      20'h0e0ed: out <= 12'h603;
      20'h0e0ee: out <= 12'h603;
      20'h0e0ef: out <= 12'h603;
      20'h0e0f0: out <= 12'h603;
      20'h0e0f1: out <= 12'h603;
      20'h0e0f2: out <= 12'h603;
      20'h0e0f3: out <= 12'h603;
      20'h0e0f4: out <= 12'h603;
      20'h0e0f5: out <= 12'h603;
      20'h0e0f6: out <= 12'h603;
      20'h0e0f7: out <= 12'h603;
      20'h0e0f8: out <= 12'h603;
      20'h0e0f9: out <= 12'h603;
      20'h0e0fa: out <= 12'h603;
      20'h0e0fb: out <= 12'h603;
      20'h0e0fc: out <= 12'h603;
      20'h0e0fd: out <= 12'h603;
      20'h0e0fe: out <= 12'h603;
      20'h0e0ff: out <= 12'h603;
      20'h0e100: out <= 12'h603;
      20'h0e101: out <= 12'h603;
      20'h0e102: out <= 12'h603;
      20'h0e103: out <= 12'h603;
      20'h0e104: out <= 12'h603;
      20'h0e105: out <= 12'h603;
      20'h0e106: out <= 12'h603;
      20'h0e107: out <= 12'h603;
      20'h0e108: out <= 12'h603;
      20'h0e109: out <= 12'h603;
      20'h0e10a: out <= 12'h603;
      20'h0e10b: out <= 12'h603;
      20'h0e10c: out <= 12'h603;
      20'h0e10d: out <= 12'h603;
      20'h0e10e: out <= 12'h603;
      20'h0e10f: out <= 12'h603;
      20'h0e110: out <= 12'hee9;
      20'h0e111: out <= 12'hf87;
      20'h0e112: out <= 12'hee9;
      20'h0e113: out <= 12'hb27;
      20'h0e114: out <= 12'hb27;
      20'h0e115: out <= 12'hb27;
      20'h0e116: out <= 12'hf87;
      20'h0e117: out <= 12'hb27;
      20'h0e118: out <= 12'h000;
      20'h0e119: out <= 12'h000;
      20'h0e11a: out <= 12'h000;
      20'h0e11b: out <= 12'h000;
      20'h0e11c: out <= 12'h000;
      20'h0e11d: out <= 12'h000;
      20'h0e11e: out <= 12'h000;
      20'h0e11f: out <= 12'h000;
      20'h0e120: out <= 12'h000;
      20'h0e121: out <= 12'h000;
      20'h0e122: out <= 12'h000;
      20'h0e123: out <= 12'h666;
      20'h0e124: out <= 12'h666;
      20'h0e125: out <= 12'hfff;
      20'h0e126: out <= 12'h666;
      20'h0e127: out <= 12'hbbb;
      20'h0e128: out <= 12'hfff;
      20'h0e129: out <= 12'hbbb;
      20'h0e12a: out <= 12'h666;
      20'h0e12b: out <= 12'h666;
      20'h0e12c: out <= 12'h666;
      20'h0e12d: out <= 12'h666;
      20'h0e12e: out <= 12'h000;
      20'h0e12f: out <= 12'h000;
      20'h0e130: out <= 12'h000;
      20'h0e131: out <= 12'h000;
      20'h0e132: out <= 12'h000;
      20'h0e133: out <= 12'h000;
      20'h0e134: out <= 12'h000;
      20'h0e135: out <= 12'h000;
      20'h0e136: out <= 12'h000;
      20'h0e137: out <= 12'h000;
      20'h0e138: out <= 12'h000;
      20'h0e139: out <= 12'h000;
      20'h0e13a: out <= 12'h000;
      20'h0e13b: out <= 12'h000;
      20'h0e13c: out <= 12'h000;
      20'h0e13d: out <= 12'h000;
      20'h0e13e: out <= 12'h000;
      20'h0e13f: out <= 12'h000;
      20'h0e140: out <= 12'h000;
      20'h0e141: out <= 12'h000;
      20'h0e142: out <= 12'h000;
      20'h0e143: out <= 12'h000;
      20'h0e144: out <= 12'h000;
      20'h0e145: out <= 12'h000;
      20'h0e146: out <= 12'h000;
      20'h0e147: out <= 12'h000;
      20'h0e148: out <= 12'h000;
      20'h0e149: out <= 12'h000;
      20'h0e14a: out <= 12'h000;
      20'h0e14b: out <= 12'h000;
      20'h0e14c: out <= 12'h000;
      20'h0e14d: out <= 12'h000;
      20'h0e14e: out <= 12'h000;
      20'h0e14f: out <= 12'h000;
      20'h0e150: out <= 12'h000;
      20'h0e151: out <= 12'h000;
      20'h0e152: out <= 12'h72f;
      20'h0e153: out <= 12'h72f;
      20'h0e154: out <= 12'h72f;
      20'h0e155: out <= 12'hc7f;
      20'h0e156: out <= 12'hc7f;
      20'h0e157: out <= 12'hc7f;
      20'h0e158: out <= 12'hc7f;
      20'h0e159: out <= 12'hc7f;
      20'h0e15a: out <= 12'hc7f;
      20'h0e15b: out <= 12'h72f;
      20'h0e15c: out <= 12'h72f;
      20'h0e15d: out <= 12'h72f;
      20'h0e15e: out <= 12'h000;
      20'h0e15f: out <= 12'h000;
      20'h0e160: out <= 12'h000;
      20'h0e161: out <= 12'h000;
      20'h0e162: out <= 12'h666;
      20'h0e163: out <= 12'h666;
      20'h0e164: out <= 12'h666;
      20'h0e165: out <= 12'hbbb;
      20'h0e166: out <= 12'hbbb;
      20'h0e167: out <= 12'hbbb;
      20'h0e168: out <= 12'hbbb;
      20'h0e169: out <= 12'hbbb;
      20'h0e16a: out <= 12'hbbb;
      20'h0e16b: out <= 12'h666;
      20'h0e16c: out <= 12'h666;
      20'h0e16d: out <= 12'h666;
      20'h0e16e: out <= 12'h000;
      20'h0e16f: out <= 12'h000;
      20'h0e170: out <= 12'h000;
      20'h0e171: out <= 12'h000;
      20'h0e172: out <= 12'h660;
      20'h0e173: out <= 12'h660;
      20'h0e174: out <= 12'h660;
      20'h0e175: out <= 12'hbb0;
      20'h0e176: out <= 12'hbb0;
      20'h0e177: out <= 12'hbb0;
      20'h0e178: out <= 12'hbb0;
      20'h0e179: out <= 12'hbb0;
      20'h0e17a: out <= 12'hbb0;
      20'h0e17b: out <= 12'h660;
      20'h0e17c: out <= 12'h660;
      20'h0e17d: out <= 12'h660;
      20'h0e17e: out <= 12'h000;
      20'h0e17f: out <= 12'h000;
      20'h0e180: out <= 12'h000;
      20'h0e181: out <= 12'h000;
      20'h0e182: out <= 12'h16d;
      20'h0e183: out <= 12'h16d;
      20'h0e184: out <= 12'h16d;
      20'h0e185: out <= 12'h6af;
      20'h0e186: out <= 12'h6af;
      20'h0e187: out <= 12'h6af;
      20'h0e188: out <= 12'h6af;
      20'h0e189: out <= 12'h6af;
      20'h0e18a: out <= 12'h6af;
      20'h0e18b: out <= 12'h16d;
      20'h0e18c: out <= 12'h16d;
      20'h0e18d: out <= 12'h16d;
      20'h0e18e: out <= 12'h000;
      20'h0e18f: out <= 12'h000;
      20'h0e190: out <= 12'h000;
      20'h0e191: out <= 12'h000;
      20'h0e192: out <= 12'h72f;
      20'h0e193: out <= 12'h72f;
      20'h0e194: out <= 12'h72f;
      20'h0e195: out <= 12'hc7f;
      20'h0e196: out <= 12'hc7f;
      20'h0e197: out <= 12'hc7f;
      20'h0e198: out <= 12'hc7f;
      20'h0e199: out <= 12'hc7f;
      20'h0e19a: out <= 12'hc7f;
      20'h0e19b: out <= 12'h72f;
      20'h0e19c: out <= 12'h72f;
      20'h0e19d: out <= 12'h72f;
      20'h0e19e: out <= 12'h000;
      20'h0e19f: out <= 12'h000;
      20'h0e1a0: out <= 12'h000;
      20'h0e1a1: out <= 12'h000;
      20'h0e1a2: out <= 12'h666;
      20'h0e1a3: out <= 12'h666;
      20'h0e1a4: out <= 12'h666;
      20'h0e1a5: out <= 12'hbbb;
      20'h0e1a6: out <= 12'hbbb;
      20'h0e1a7: out <= 12'hbbb;
      20'h0e1a8: out <= 12'hbbb;
      20'h0e1a9: out <= 12'hbbb;
      20'h0e1aa: out <= 12'hbbb;
      20'h0e1ab: out <= 12'h666;
      20'h0e1ac: out <= 12'h666;
      20'h0e1ad: out <= 12'h666;
      20'h0e1ae: out <= 12'h000;
      20'h0e1af: out <= 12'h000;
      20'h0e1b0: out <= 12'h000;
      20'h0e1b1: out <= 12'h000;
      20'h0e1b2: out <= 12'h16d;
      20'h0e1b3: out <= 12'h16d;
      20'h0e1b4: out <= 12'h16d;
      20'h0e1b5: out <= 12'h6af;
      20'h0e1b6: out <= 12'h6af;
      20'h0e1b7: out <= 12'h6af;
      20'h0e1b8: out <= 12'h6af;
      20'h0e1b9: out <= 12'h6af;
      20'h0e1ba: out <= 12'h6af;
      20'h0e1bb: out <= 12'h16d;
      20'h0e1bc: out <= 12'h16d;
      20'h0e1bd: out <= 12'h16d;
      20'h0e1be: out <= 12'h000;
      20'h0e1bf: out <= 12'h000;
      20'h0e1c0: out <= 12'h000;
      20'h0e1c1: out <= 12'h000;
      20'h0e1c2: out <= 12'h660;
      20'h0e1c3: out <= 12'h660;
      20'h0e1c4: out <= 12'h660;
      20'h0e1c5: out <= 12'hbb0;
      20'h0e1c6: out <= 12'hbb0;
      20'h0e1c7: out <= 12'hbb0;
      20'h0e1c8: out <= 12'hbb0;
      20'h0e1c9: out <= 12'hbb0;
      20'h0e1ca: out <= 12'hbb0;
      20'h0e1cb: out <= 12'h660;
      20'h0e1cc: out <= 12'h660;
      20'h0e1cd: out <= 12'h660;
      20'h0e1ce: out <= 12'h000;
      20'h0e1cf: out <= 12'h000;
      20'h0e1d0: out <= 12'h603;
      20'h0e1d1: out <= 12'h603;
      20'h0e1d2: out <= 12'h603;
      20'h0e1d3: out <= 12'h603;
      20'h0e1d4: out <= 12'h603;
      20'h0e1d5: out <= 12'h603;
      20'h0e1d6: out <= 12'h603;
      20'h0e1d7: out <= 12'h603;
      20'h0e1d8: out <= 12'h603;
      20'h0e1d9: out <= 12'h603;
      20'h0e1da: out <= 12'h603;
      20'h0e1db: out <= 12'h603;
      20'h0e1dc: out <= 12'h603;
      20'h0e1dd: out <= 12'h603;
      20'h0e1de: out <= 12'h603;
      20'h0e1df: out <= 12'h603;
      20'h0e1e0: out <= 12'h603;
      20'h0e1e1: out <= 12'h603;
      20'h0e1e2: out <= 12'h603;
      20'h0e1e3: out <= 12'h603;
      20'h0e1e4: out <= 12'h603;
      20'h0e1e5: out <= 12'h603;
      20'h0e1e6: out <= 12'h603;
      20'h0e1e7: out <= 12'h603;
      20'h0e1e8: out <= 12'h603;
      20'h0e1e9: out <= 12'h603;
      20'h0e1ea: out <= 12'h603;
      20'h0e1eb: out <= 12'h603;
      20'h0e1ec: out <= 12'h603;
      20'h0e1ed: out <= 12'h603;
      20'h0e1ee: out <= 12'h603;
      20'h0e1ef: out <= 12'h603;
      20'h0e1f0: out <= 12'h603;
      20'h0e1f1: out <= 12'h603;
      20'h0e1f2: out <= 12'h603;
      20'h0e1f3: out <= 12'h603;
      20'h0e1f4: out <= 12'h603;
      20'h0e1f5: out <= 12'h603;
      20'h0e1f6: out <= 12'h603;
      20'h0e1f7: out <= 12'h603;
      20'h0e1f8: out <= 12'h603;
      20'h0e1f9: out <= 12'h603;
      20'h0e1fa: out <= 12'h603;
      20'h0e1fb: out <= 12'h603;
      20'h0e1fc: out <= 12'h603;
      20'h0e1fd: out <= 12'h603;
      20'h0e1fe: out <= 12'h603;
      20'h0e1ff: out <= 12'h603;
      20'h0e200: out <= 12'h603;
      20'h0e201: out <= 12'h603;
      20'h0e202: out <= 12'h603;
      20'h0e203: out <= 12'h603;
      20'h0e204: out <= 12'h603;
      20'h0e205: out <= 12'h603;
      20'h0e206: out <= 12'h603;
      20'h0e207: out <= 12'h603;
      20'h0e208: out <= 12'h603;
      20'h0e209: out <= 12'h603;
      20'h0e20a: out <= 12'h603;
      20'h0e20b: out <= 12'h603;
      20'h0e20c: out <= 12'h603;
      20'h0e20d: out <= 12'h603;
      20'h0e20e: out <= 12'h603;
      20'h0e20f: out <= 12'h603;
      20'h0e210: out <= 12'h603;
      20'h0e211: out <= 12'h603;
      20'h0e212: out <= 12'h603;
      20'h0e213: out <= 12'h603;
      20'h0e214: out <= 12'h603;
      20'h0e215: out <= 12'h603;
      20'h0e216: out <= 12'h603;
      20'h0e217: out <= 12'h603;
      20'h0e218: out <= 12'h603;
      20'h0e219: out <= 12'h603;
      20'h0e21a: out <= 12'h603;
      20'h0e21b: out <= 12'h603;
      20'h0e21c: out <= 12'h603;
      20'h0e21d: out <= 12'h603;
      20'h0e21e: out <= 12'h603;
      20'h0e21f: out <= 12'h603;
      20'h0e220: out <= 12'h603;
      20'h0e221: out <= 12'h603;
      20'h0e222: out <= 12'h603;
      20'h0e223: out <= 12'h603;
      20'h0e224: out <= 12'h603;
      20'h0e225: out <= 12'h603;
      20'h0e226: out <= 12'h603;
      20'h0e227: out <= 12'h603;
      20'h0e228: out <= 12'hee9;
      20'h0e229: out <= 12'hf87;
      20'h0e22a: out <= 12'hf87;
      20'h0e22b: out <= 12'hf87;
      20'h0e22c: out <= 12'hf87;
      20'h0e22d: out <= 12'hf87;
      20'h0e22e: out <= 12'hf87;
      20'h0e22f: out <= 12'hb27;
      20'h0e230: out <= 12'h000;
      20'h0e231: out <= 12'h000;
      20'h0e232: out <= 12'h000;
      20'h0e233: out <= 12'h000;
      20'h0e234: out <= 12'h000;
      20'h0e235: out <= 12'h000;
      20'h0e236: out <= 12'h000;
      20'h0e237: out <= 12'h000;
      20'h0e238: out <= 12'h000;
      20'h0e239: out <= 12'h000;
      20'h0e23a: out <= 12'h666;
      20'h0e23b: out <= 12'hbbb;
      20'h0e23c: out <= 12'h666;
      20'h0e23d: out <= 12'hfff;
      20'h0e23e: out <= 12'h666;
      20'h0e23f: out <= 12'hbbb;
      20'h0e240: out <= 12'hfff;
      20'h0e241: out <= 12'hbbb;
      20'h0e242: out <= 12'h666;
      20'h0e243: out <= 12'h666;
      20'h0e244: out <= 12'h666;
      20'h0e245: out <= 12'hbbb;
      20'h0e246: out <= 12'h666;
      20'h0e247: out <= 12'h000;
      20'h0e248: out <= 12'h000;
      20'h0e249: out <= 12'h000;
      20'h0e24a: out <= 12'h000;
      20'h0e24b: out <= 12'h000;
      20'h0e24c: out <= 12'h000;
      20'h0e24d: out <= 12'h000;
      20'h0e24e: out <= 12'h000;
      20'h0e24f: out <= 12'h000;
      20'h0e250: out <= 12'h000;
      20'h0e251: out <= 12'h000;
      20'h0e252: out <= 12'h000;
      20'h0e253: out <= 12'h000;
      20'h0e254: out <= 12'h000;
      20'h0e255: out <= 12'h000;
      20'h0e256: out <= 12'h000;
      20'h0e257: out <= 12'h000;
      20'h0e258: out <= 12'h000;
      20'h0e259: out <= 12'h000;
      20'h0e25a: out <= 12'h000;
      20'h0e25b: out <= 12'h000;
      20'h0e25c: out <= 12'h000;
      20'h0e25d: out <= 12'h000;
      20'h0e25e: out <= 12'h000;
      20'h0e25f: out <= 12'h000;
      20'h0e260: out <= 12'h000;
      20'h0e261: out <= 12'h000;
      20'h0e262: out <= 12'h000;
      20'h0e263: out <= 12'h000;
      20'h0e264: out <= 12'h000;
      20'h0e265: out <= 12'h000;
      20'h0e266: out <= 12'h000;
      20'h0e267: out <= 12'h000;
      20'h0e268: out <= 12'h000;
      20'h0e269: out <= 12'h000;
      20'h0e26a: out <= 12'h000;
      20'h0e26b: out <= 12'h000;
      20'h0e26c: out <= 12'h000;
      20'h0e26d: out <= 12'h000;
      20'h0e26e: out <= 12'h000;
      20'h0e26f: out <= 12'h000;
      20'h0e270: out <= 12'h000;
      20'h0e271: out <= 12'h000;
      20'h0e272: out <= 12'h000;
      20'h0e273: out <= 12'h000;
      20'h0e274: out <= 12'h000;
      20'h0e275: out <= 12'h000;
      20'h0e276: out <= 12'h000;
      20'h0e277: out <= 12'h000;
      20'h0e278: out <= 12'h000;
      20'h0e279: out <= 12'h000;
      20'h0e27a: out <= 12'h000;
      20'h0e27b: out <= 12'h000;
      20'h0e27c: out <= 12'h000;
      20'h0e27d: out <= 12'h000;
      20'h0e27e: out <= 12'h000;
      20'h0e27f: out <= 12'h000;
      20'h0e280: out <= 12'h000;
      20'h0e281: out <= 12'h000;
      20'h0e282: out <= 12'h000;
      20'h0e283: out <= 12'h000;
      20'h0e284: out <= 12'h000;
      20'h0e285: out <= 12'h000;
      20'h0e286: out <= 12'h000;
      20'h0e287: out <= 12'h000;
      20'h0e288: out <= 12'h000;
      20'h0e289: out <= 12'h000;
      20'h0e28a: out <= 12'h000;
      20'h0e28b: out <= 12'h000;
      20'h0e28c: out <= 12'h000;
      20'h0e28d: out <= 12'h000;
      20'h0e28e: out <= 12'h000;
      20'h0e28f: out <= 12'h000;
      20'h0e290: out <= 12'h000;
      20'h0e291: out <= 12'h000;
      20'h0e292: out <= 12'h000;
      20'h0e293: out <= 12'h000;
      20'h0e294: out <= 12'h000;
      20'h0e295: out <= 12'h000;
      20'h0e296: out <= 12'h000;
      20'h0e297: out <= 12'h000;
      20'h0e298: out <= 12'h000;
      20'h0e299: out <= 12'h000;
      20'h0e29a: out <= 12'h000;
      20'h0e29b: out <= 12'h000;
      20'h0e29c: out <= 12'h000;
      20'h0e29d: out <= 12'h000;
      20'h0e29e: out <= 12'h000;
      20'h0e29f: out <= 12'h000;
      20'h0e2a0: out <= 12'h000;
      20'h0e2a1: out <= 12'h000;
      20'h0e2a2: out <= 12'h000;
      20'h0e2a3: out <= 12'h000;
      20'h0e2a4: out <= 12'h000;
      20'h0e2a5: out <= 12'h000;
      20'h0e2a6: out <= 12'h000;
      20'h0e2a7: out <= 12'h000;
      20'h0e2a8: out <= 12'h000;
      20'h0e2a9: out <= 12'h000;
      20'h0e2aa: out <= 12'h000;
      20'h0e2ab: out <= 12'h000;
      20'h0e2ac: out <= 12'h000;
      20'h0e2ad: out <= 12'h000;
      20'h0e2ae: out <= 12'h000;
      20'h0e2af: out <= 12'h000;
      20'h0e2b0: out <= 12'h000;
      20'h0e2b1: out <= 12'h000;
      20'h0e2b2: out <= 12'h000;
      20'h0e2b3: out <= 12'h000;
      20'h0e2b4: out <= 12'h000;
      20'h0e2b5: out <= 12'h000;
      20'h0e2b6: out <= 12'h000;
      20'h0e2b7: out <= 12'h000;
      20'h0e2b8: out <= 12'h000;
      20'h0e2b9: out <= 12'h000;
      20'h0e2ba: out <= 12'h000;
      20'h0e2bb: out <= 12'h000;
      20'h0e2bc: out <= 12'h000;
      20'h0e2bd: out <= 12'h000;
      20'h0e2be: out <= 12'h000;
      20'h0e2bf: out <= 12'h000;
      20'h0e2c0: out <= 12'h000;
      20'h0e2c1: out <= 12'h000;
      20'h0e2c2: out <= 12'h000;
      20'h0e2c3: out <= 12'h000;
      20'h0e2c4: out <= 12'h000;
      20'h0e2c5: out <= 12'h000;
      20'h0e2c6: out <= 12'h000;
      20'h0e2c7: out <= 12'h000;
      20'h0e2c8: out <= 12'h000;
      20'h0e2c9: out <= 12'h000;
      20'h0e2ca: out <= 12'h000;
      20'h0e2cb: out <= 12'h000;
      20'h0e2cc: out <= 12'h000;
      20'h0e2cd: out <= 12'h000;
      20'h0e2ce: out <= 12'h000;
      20'h0e2cf: out <= 12'h000;
      20'h0e2d0: out <= 12'h000;
      20'h0e2d1: out <= 12'h000;
      20'h0e2d2: out <= 12'h000;
      20'h0e2d3: out <= 12'h000;
      20'h0e2d4: out <= 12'h000;
      20'h0e2d5: out <= 12'h000;
      20'h0e2d6: out <= 12'h000;
      20'h0e2d7: out <= 12'h000;
      20'h0e2d8: out <= 12'h000;
      20'h0e2d9: out <= 12'h000;
      20'h0e2da: out <= 12'h000;
      20'h0e2db: out <= 12'h000;
      20'h0e2dc: out <= 12'h000;
      20'h0e2dd: out <= 12'h000;
      20'h0e2de: out <= 12'h000;
      20'h0e2df: out <= 12'h000;
      20'h0e2e0: out <= 12'h000;
      20'h0e2e1: out <= 12'h000;
      20'h0e2e2: out <= 12'h000;
      20'h0e2e3: out <= 12'h000;
      20'h0e2e4: out <= 12'h000;
      20'h0e2e5: out <= 12'h000;
      20'h0e2e6: out <= 12'h000;
      20'h0e2e7: out <= 12'h000;
      20'h0e2e8: out <= 12'h603;
      20'h0e2e9: out <= 12'h603;
      20'h0e2ea: out <= 12'h603;
      20'h0e2eb: out <= 12'h603;
      20'h0e2ec: out <= 12'h603;
      20'h0e2ed: out <= 12'h603;
      20'h0e2ee: out <= 12'h603;
      20'h0e2ef: out <= 12'h603;
      20'h0e2f0: out <= 12'h603;
      20'h0e2f1: out <= 12'h603;
      20'h0e2f2: out <= 12'h603;
      20'h0e2f3: out <= 12'h603;
      20'h0e2f4: out <= 12'h603;
      20'h0e2f5: out <= 12'h603;
      20'h0e2f6: out <= 12'h603;
      20'h0e2f7: out <= 12'h603;
      20'h0e2f8: out <= 12'h603;
      20'h0e2f9: out <= 12'h603;
      20'h0e2fa: out <= 12'h603;
      20'h0e2fb: out <= 12'h603;
      20'h0e2fc: out <= 12'h603;
      20'h0e2fd: out <= 12'h603;
      20'h0e2fe: out <= 12'h603;
      20'h0e2ff: out <= 12'h603;
      20'h0e300: out <= 12'h603;
      20'h0e301: out <= 12'h603;
      20'h0e302: out <= 12'h603;
      20'h0e303: out <= 12'h603;
      20'h0e304: out <= 12'h603;
      20'h0e305: out <= 12'h603;
      20'h0e306: out <= 12'h603;
      20'h0e307: out <= 12'h603;
      20'h0e308: out <= 12'h603;
      20'h0e309: out <= 12'h603;
      20'h0e30a: out <= 12'h603;
      20'h0e30b: out <= 12'h603;
      20'h0e30c: out <= 12'h603;
      20'h0e30d: out <= 12'h603;
      20'h0e30e: out <= 12'h603;
      20'h0e30f: out <= 12'h603;
      20'h0e310: out <= 12'h603;
      20'h0e311: out <= 12'h603;
      20'h0e312: out <= 12'h603;
      20'h0e313: out <= 12'h603;
      20'h0e314: out <= 12'h603;
      20'h0e315: out <= 12'h603;
      20'h0e316: out <= 12'h603;
      20'h0e317: out <= 12'h603;
      20'h0e318: out <= 12'h603;
      20'h0e319: out <= 12'h603;
      20'h0e31a: out <= 12'h603;
      20'h0e31b: out <= 12'h603;
      20'h0e31c: out <= 12'h603;
      20'h0e31d: out <= 12'h603;
      20'h0e31e: out <= 12'h603;
      20'h0e31f: out <= 12'h603;
      20'h0e320: out <= 12'h603;
      20'h0e321: out <= 12'h603;
      20'h0e322: out <= 12'h603;
      20'h0e323: out <= 12'h603;
      20'h0e324: out <= 12'h603;
      20'h0e325: out <= 12'h603;
      20'h0e326: out <= 12'h603;
      20'h0e327: out <= 12'h603;
      20'h0e328: out <= 12'h603;
      20'h0e329: out <= 12'h603;
      20'h0e32a: out <= 12'h603;
      20'h0e32b: out <= 12'h603;
      20'h0e32c: out <= 12'h603;
      20'h0e32d: out <= 12'h603;
      20'h0e32e: out <= 12'h603;
      20'h0e32f: out <= 12'h603;
      20'h0e330: out <= 12'h603;
      20'h0e331: out <= 12'h603;
      20'h0e332: out <= 12'h603;
      20'h0e333: out <= 12'h603;
      20'h0e334: out <= 12'h603;
      20'h0e335: out <= 12'h603;
      20'h0e336: out <= 12'h603;
      20'h0e337: out <= 12'h603;
      20'h0e338: out <= 12'h603;
      20'h0e339: out <= 12'h603;
      20'h0e33a: out <= 12'h603;
      20'h0e33b: out <= 12'h603;
      20'h0e33c: out <= 12'h603;
      20'h0e33d: out <= 12'h603;
      20'h0e33e: out <= 12'h603;
      20'h0e33f: out <= 12'h603;
      20'h0e340: out <= 12'hb27;
      20'h0e341: out <= 12'hb27;
      20'h0e342: out <= 12'hb27;
      20'h0e343: out <= 12'hb27;
      20'h0e344: out <= 12'hb27;
      20'h0e345: out <= 12'hb27;
      20'h0e346: out <= 12'hb27;
      20'h0e347: out <= 12'hb27;
      20'h0e348: out <= 12'h000;
      20'h0e349: out <= 12'h000;
      20'h0e34a: out <= 12'h000;
      20'h0e34b: out <= 12'h000;
      20'h0e34c: out <= 12'h000;
      20'h0e34d: out <= 12'h000;
      20'h0e34e: out <= 12'h000;
      20'h0e34f: out <= 12'h000;
      20'h0e350: out <= 12'h000;
      20'h0e351: out <= 12'h000;
      20'h0e352: out <= 12'h000;
      20'h0e353: out <= 12'h666;
      20'h0e354: out <= 12'h666;
      20'h0e355: out <= 12'hfff;
      20'h0e356: out <= 12'hbbb;
      20'h0e357: out <= 12'h666;
      20'h0e358: out <= 12'h666;
      20'h0e359: out <= 12'h666;
      20'h0e35a: out <= 12'h666;
      20'h0e35b: out <= 12'h666;
      20'h0e35c: out <= 12'h666;
      20'h0e35d: out <= 12'h666;
      20'h0e35e: out <= 12'h000;
      20'h0e35f: out <= 12'h000;
      20'h0e360: out <= 12'h000;
      20'h0e361: out <= 12'h000;
      20'h0e362: out <= 12'h000;
      20'h0e363: out <= 12'h000;
      20'h0e364: out <= 12'h000;
      20'h0e365: out <= 12'h000;
      20'h0e366: out <= 12'h000;
      20'h0e367: out <= 12'h000;
      20'h0e368: out <= 12'h000;
      20'h0e369: out <= 12'h000;
      20'h0e36a: out <= 12'h000;
      20'h0e36b: out <= 12'h000;
      20'h0e36c: out <= 12'h000;
      20'h0e36d: out <= 12'h000;
      20'h0e36e: out <= 12'h000;
      20'h0e36f: out <= 12'h000;
      20'h0e370: out <= 12'h000;
      20'h0e371: out <= 12'h000;
      20'h0e372: out <= 12'h000;
      20'h0e373: out <= 12'h000;
      20'h0e374: out <= 12'h000;
      20'h0e375: out <= 12'h000;
      20'h0e376: out <= 12'h000;
      20'h0e377: out <= 12'h000;
      20'h0e378: out <= 12'h000;
      20'h0e379: out <= 12'h000;
      20'h0e37a: out <= 12'h000;
      20'h0e37b: out <= 12'h000;
      20'h0e37c: out <= 12'h000;
      20'h0e37d: out <= 12'h000;
      20'h0e37e: out <= 12'h000;
      20'h0e37f: out <= 12'h000;
      20'h0e380: out <= 12'hfff;
      20'h0e381: out <= 12'hfff;
      20'h0e382: out <= 12'hfff;
      20'h0e383: out <= 12'hfff;
      20'h0e384: out <= 12'hfff;
      20'h0e385: out <= 12'hfff;
      20'h0e386: out <= 12'hfff;
      20'h0e387: out <= 12'hfff;
      20'h0e388: out <= 12'hfff;
      20'h0e389: out <= 12'hfff;
      20'h0e38a: out <= 12'hfff;
      20'h0e38b: out <= 12'hfff;
      20'h0e38c: out <= 12'hfff;
      20'h0e38d: out <= 12'hfff;
      20'h0e38e: out <= 12'hfff;
      20'h0e38f: out <= 12'hfff;
      20'h0e390: out <= 12'hfff;
      20'h0e391: out <= 12'hfff;
      20'h0e392: out <= 12'hfff;
      20'h0e393: out <= 12'hfff;
      20'h0e394: out <= 12'hfff;
      20'h0e395: out <= 12'hfff;
      20'h0e396: out <= 12'hfff;
      20'h0e397: out <= 12'hfff;
      20'h0e398: out <= 12'hfff;
      20'h0e399: out <= 12'hfff;
      20'h0e39a: out <= 12'hfff;
      20'h0e39b: out <= 12'hfff;
      20'h0e39c: out <= 12'hfff;
      20'h0e39d: out <= 12'hfff;
      20'h0e39e: out <= 12'hfff;
      20'h0e39f: out <= 12'hfff;
      20'h0e3a0: out <= 12'hfff;
      20'h0e3a1: out <= 12'hfff;
      20'h0e3a2: out <= 12'hfff;
      20'h0e3a3: out <= 12'hfff;
      20'h0e3a4: out <= 12'hfff;
      20'h0e3a5: out <= 12'hfff;
      20'h0e3a6: out <= 12'hfff;
      20'h0e3a7: out <= 12'hfff;
      20'h0e3a8: out <= 12'hfff;
      20'h0e3a9: out <= 12'hfff;
      20'h0e3aa: out <= 12'hfff;
      20'h0e3ab: out <= 12'hfff;
      20'h0e3ac: out <= 12'hfff;
      20'h0e3ad: out <= 12'hfff;
      20'h0e3ae: out <= 12'hfff;
      20'h0e3af: out <= 12'hfff;
      20'h0e3b0: out <= 12'h603;
      20'h0e3b1: out <= 12'h603;
      20'h0e3b2: out <= 12'h603;
      20'h0e3b3: out <= 12'h603;
      20'h0e3b4: out <= 12'h603;
      20'h0e3b5: out <= 12'h603;
      20'h0e3b6: out <= 12'h603;
      20'h0e3b7: out <= 12'h603;
      20'h0e3b8: out <= 12'h603;
      20'h0e3b9: out <= 12'h603;
      20'h0e3ba: out <= 12'h603;
      20'h0e3bb: out <= 12'h603;
      20'h0e3bc: out <= 12'h603;
      20'h0e3bd: out <= 12'h603;
      20'h0e3be: out <= 12'h603;
      20'h0e3bf: out <= 12'h603;
      20'h0e3c0: out <= 12'h603;
      20'h0e3c1: out <= 12'h603;
      20'h0e3c2: out <= 12'h603;
      20'h0e3c3: out <= 12'h603;
      20'h0e3c4: out <= 12'h603;
      20'h0e3c5: out <= 12'h603;
      20'h0e3c6: out <= 12'h603;
      20'h0e3c7: out <= 12'h603;
      20'h0e3c8: out <= 12'h603;
      20'h0e3c9: out <= 12'h603;
      20'h0e3ca: out <= 12'h603;
      20'h0e3cb: out <= 12'h603;
      20'h0e3cc: out <= 12'h603;
      20'h0e3cd: out <= 12'h603;
      20'h0e3ce: out <= 12'h603;
      20'h0e3cf: out <= 12'h603;
      20'h0e3d0: out <= 12'h603;
      20'h0e3d1: out <= 12'h603;
      20'h0e3d2: out <= 12'h603;
      20'h0e3d3: out <= 12'h603;
      20'h0e3d4: out <= 12'h603;
      20'h0e3d5: out <= 12'h603;
      20'h0e3d6: out <= 12'h603;
      20'h0e3d7: out <= 12'h603;
      20'h0e3d8: out <= 12'hfff;
      20'h0e3d9: out <= 12'hfff;
      20'h0e3da: out <= 12'hfff;
      20'h0e3db: out <= 12'hfff;
      20'h0e3dc: out <= 12'hfff;
      20'h0e3dd: out <= 12'hfff;
      20'h0e3de: out <= 12'hfff;
      20'h0e3df: out <= 12'hfff;
      20'h0e3e0: out <= 12'hfff;
      20'h0e3e1: out <= 12'hfff;
      20'h0e3e2: out <= 12'hfff;
      20'h0e3e3: out <= 12'hfff;
      20'h0e3e4: out <= 12'hfff;
      20'h0e3e5: out <= 12'hfff;
      20'h0e3e6: out <= 12'hfff;
      20'h0e3e7: out <= 12'hfff;
      20'h0e3e8: out <= 12'hfff;
      20'h0e3e9: out <= 12'hfff;
      20'h0e3ea: out <= 12'hfff;
      20'h0e3eb: out <= 12'hfff;
      20'h0e3ec: out <= 12'hfff;
      20'h0e3ed: out <= 12'hfff;
      20'h0e3ee: out <= 12'hfff;
      20'h0e3ef: out <= 12'hfff;
      20'h0e3f0: out <= 12'hfff;
      20'h0e3f1: out <= 12'hfff;
      20'h0e3f2: out <= 12'hfff;
      20'h0e3f3: out <= 12'hfff;
      20'h0e3f4: out <= 12'hfff;
      20'h0e3f5: out <= 12'hfff;
      20'h0e3f6: out <= 12'hfff;
      20'h0e3f7: out <= 12'hfff;
      20'h0e3f8: out <= 12'hfff;
      20'h0e3f9: out <= 12'hfff;
      20'h0e3fa: out <= 12'hfff;
      20'h0e3fb: out <= 12'hfff;
      20'h0e3fc: out <= 12'hfff;
      20'h0e3fd: out <= 12'hfff;
      20'h0e3fe: out <= 12'hfff;
      20'h0e3ff: out <= 12'h72f;
      20'h0e400: out <= 12'h603;
      20'h0e401: out <= 12'h603;
      20'h0e402: out <= 12'h603;
      20'h0e403: out <= 12'h603;
      20'h0e404: out <= 12'h603;
      20'h0e405: out <= 12'h603;
      20'h0e406: out <= 12'h603;
      20'h0e407: out <= 12'h603;
      20'h0e408: out <= 12'h603;
      20'h0e409: out <= 12'h603;
      20'h0e40a: out <= 12'h603;
      20'h0e40b: out <= 12'h603;
      20'h0e40c: out <= 12'h603;
      20'h0e40d: out <= 12'h603;
      20'h0e40e: out <= 12'h603;
      20'h0e40f: out <= 12'h603;
      20'h0e410: out <= 12'h603;
      20'h0e411: out <= 12'h603;
      20'h0e412: out <= 12'h603;
      20'h0e413: out <= 12'h603;
      20'h0e414: out <= 12'h603;
      20'h0e415: out <= 12'h603;
      20'h0e416: out <= 12'h603;
      20'h0e417: out <= 12'h603;
      20'h0e418: out <= 12'h603;
      20'h0e419: out <= 12'h603;
      20'h0e41a: out <= 12'h603;
      20'h0e41b: out <= 12'h603;
      20'h0e41c: out <= 12'h603;
      20'h0e41d: out <= 12'h603;
      20'h0e41e: out <= 12'h603;
      20'h0e41f: out <= 12'h603;
      20'h0e420: out <= 12'h603;
      20'h0e421: out <= 12'h603;
      20'h0e422: out <= 12'h603;
      20'h0e423: out <= 12'h603;
      20'h0e424: out <= 12'h603;
      20'h0e425: out <= 12'h603;
      20'h0e426: out <= 12'h603;
      20'h0e427: out <= 12'h603;
      20'h0e428: out <= 12'h603;
      20'h0e429: out <= 12'h603;
      20'h0e42a: out <= 12'h603;
      20'h0e42b: out <= 12'h603;
      20'h0e42c: out <= 12'h603;
      20'h0e42d: out <= 12'h603;
      20'h0e42e: out <= 12'h603;
      20'h0e42f: out <= 12'h603;
      20'h0e430: out <= 12'h603;
      20'h0e431: out <= 12'h603;
      20'h0e432: out <= 12'h603;
      20'h0e433: out <= 12'h603;
      20'h0e434: out <= 12'h603;
      20'h0e435: out <= 12'h603;
      20'h0e436: out <= 12'h603;
      20'h0e437: out <= 12'h603;
      20'h0e438: out <= 12'h603;
      20'h0e439: out <= 12'h603;
      20'h0e43a: out <= 12'h603;
      20'h0e43b: out <= 12'h603;
      20'h0e43c: out <= 12'h603;
      20'h0e43d: out <= 12'h603;
      20'h0e43e: out <= 12'h603;
      20'h0e43f: out <= 12'h603;
      20'h0e440: out <= 12'h603;
      20'h0e441: out <= 12'h603;
      20'h0e442: out <= 12'h603;
      20'h0e443: out <= 12'h603;
      20'h0e444: out <= 12'h603;
      20'h0e445: out <= 12'h603;
      20'h0e446: out <= 12'h603;
      20'h0e447: out <= 12'h603;
      20'h0e448: out <= 12'h603;
      20'h0e449: out <= 12'h603;
      20'h0e44a: out <= 12'h603;
      20'h0e44b: out <= 12'h603;
      20'h0e44c: out <= 12'h603;
      20'h0e44d: out <= 12'h603;
      20'h0e44e: out <= 12'h603;
      20'h0e44f: out <= 12'h603;
      20'h0e450: out <= 12'h603;
      20'h0e451: out <= 12'h603;
      20'h0e452: out <= 12'h603;
      20'h0e453: out <= 12'h603;
      20'h0e454: out <= 12'h603;
      20'h0e455: out <= 12'h603;
      20'h0e456: out <= 12'h603;
      20'h0e457: out <= 12'h603;
      20'h0e458: out <= 12'hee9;
      20'h0e459: out <= 12'hee9;
      20'h0e45a: out <= 12'hee9;
      20'h0e45b: out <= 12'hee9;
      20'h0e45c: out <= 12'hee9;
      20'h0e45d: out <= 12'hee9;
      20'h0e45e: out <= 12'hee9;
      20'h0e45f: out <= 12'hb27;
      20'h0e460: out <= 12'h000;
      20'h0e461: out <= 12'h000;
      20'h0e462: out <= 12'h000;
      20'h0e463: out <= 12'h000;
      20'h0e464: out <= 12'h000;
      20'h0e465: out <= 12'h000;
      20'h0e466: out <= 12'h000;
      20'h0e467: out <= 12'h000;
      20'h0e468: out <= 12'h000;
      20'h0e469: out <= 12'h000;
      20'h0e46a: out <= 12'h666;
      20'h0e46b: out <= 12'hbbb;
      20'h0e46c: out <= 12'h666;
      20'h0e46d: out <= 12'hfff;
      20'h0e46e: out <= 12'h666;
      20'h0e46f: out <= 12'hfff;
      20'h0e470: out <= 12'hfff;
      20'h0e471: out <= 12'hbbb;
      20'h0e472: out <= 12'h666;
      20'h0e473: out <= 12'h666;
      20'h0e474: out <= 12'h666;
      20'h0e475: out <= 12'hbbb;
      20'h0e476: out <= 12'h666;
      20'h0e477: out <= 12'h000;
      20'h0e478: out <= 12'h000;
      20'h0e479: out <= 12'h000;
      20'h0e47a: out <= 12'h000;
      20'h0e47b: out <= 12'h000;
      20'h0e47c: out <= 12'h000;
      20'h0e47d: out <= 12'h000;
      20'h0e47e: out <= 12'h000;
      20'h0e47f: out <= 12'h000;
      20'h0e480: out <= 12'h999;
      20'h0e481: out <= 12'h999;
      20'h0e482: out <= 12'h999;
      20'h0e483: out <= 12'h999;
      20'h0e484: out <= 12'h999;
      20'h0e485: out <= 12'h999;
      20'h0e486: out <= 12'h999;
      20'h0e487: out <= 12'h999;
      20'h0e488: out <= 12'hbbb;
      20'h0e489: out <= 12'hbbb;
      20'h0e48a: out <= 12'hbbb;
      20'h0e48b: out <= 12'hbbb;
      20'h0e48c: out <= 12'hbbb;
      20'h0e48d: out <= 12'hbbb;
      20'h0e48e: out <= 12'hbbb;
      20'h0e48f: out <= 12'hbbb;
      20'h0e490: out <= 12'h000;
      20'h0e491: out <= 12'h000;
      20'h0e492: out <= 12'h000;
      20'h0e493: out <= 12'h000;
      20'h0e494: out <= 12'h000;
      20'h0e495: out <= 12'h000;
      20'h0e496: out <= 12'h000;
      20'h0e497: out <= 12'h000;
      20'h0e498: out <= 12'hfff;
      20'h0e499: out <= 12'hfff;
      20'h0e49a: out <= 12'hfff;
      20'h0e49b: out <= 12'hfff;
      20'h0e49c: out <= 12'hfff;
      20'h0e49d: out <= 12'hfff;
      20'h0e49e: out <= 12'hfff;
      20'h0e49f: out <= 12'hfff;
      20'h0e4a0: out <= 12'hfff;
      20'h0e4a1: out <= 12'hfff;
      20'h0e4a2: out <= 12'hfff;
      20'h0e4a3: out <= 12'hfff;
      20'h0e4a4: out <= 12'hfff;
      20'h0e4a5: out <= 12'hfff;
      20'h0e4a6: out <= 12'hfff;
      20'h0e4a7: out <= 12'hfff;
      20'h0e4a8: out <= 12'hfff;
      20'h0e4a9: out <= 12'hfff;
      20'h0e4aa: out <= 12'hfff;
      20'h0e4ab: out <= 12'hfff;
      20'h0e4ac: out <= 12'hfff;
      20'h0e4ad: out <= 12'hfff;
      20'h0e4ae: out <= 12'hfff;
      20'h0e4af: out <= 12'hfff;
      20'h0e4b0: out <= 12'hfff;
      20'h0e4b1: out <= 12'hfff;
      20'h0e4b2: out <= 12'hfff;
      20'h0e4b3: out <= 12'hfff;
      20'h0e4b4: out <= 12'hfff;
      20'h0e4b5: out <= 12'hfff;
      20'h0e4b6: out <= 12'hfff;
      20'h0e4b7: out <= 12'hfff;
      20'h0e4b8: out <= 12'hfff;
      20'h0e4b9: out <= 12'hfff;
      20'h0e4ba: out <= 12'hfff;
      20'h0e4bb: out <= 12'hfff;
      20'h0e4bc: out <= 12'hfff;
      20'h0e4bd: out <= 12'hfff;
      20'h0e4be: out <= 12'hfff;
      20'h0e4bf: out <= 12'hfff;
      20'h0e4c0: out <= 12'hfff;
      20'h0e4c1: out <= 12'hfff;
      20'h0e4c2: out <= 12'hfff;
      20'h0e4c3: out <= 12'hfff;
      20'h0e4c4: out <= 12'hfff;
      20'h0e4c5: out <= 12'hfff;
      20'h0e4c6: out <= 12'hfff;
      20'h0e4c7: out <= 12'h666;
      20'h0e4c8: out <= 12'h603;
      20'h0e4c9: out <= 12'h603;
      20'h0e4ca: out <= 12'h603;
      20'h0e4cb: out <= 12'h603;
      20'h0e4cc: out <= 12'h603;
      20'h0e4cd: out <= 12'h603;
      20'h0e4ce: out <= 12'h603;
      20'h0e4cf: out <= 12'h603;
      20'h0e4d0: out <= 12'h603;
      20'h0e4d1: out <= 12'h603;
      20'h0e4d2: out <= 12'h603;
      20'h0e4d3: out <= 12'h603;
      20'h0e4d4: out <= 12'h603;
      20'h0e4d5: out <= 12'h603;
      20'h0e4d6: out <= 12'h603;
      20'h0e4d7: out <= 12'h603;
      20'h0e4d8: out <= 12'h603;
      20'h0e4d9: out <= 12'h603;
      20'h0e4da: out <= 12'h603;
      20'h0e4db: out <= 12'h603;
      20'h0e4dc: out <= 12'h603;
      20'h0e4dd: out <= 12'h603;
      20'h0e4de: out <= 12'h603;
      20'h0e4df: out <= 12'h603;
      20'h0e4e0: out <= 12'h603;
      20'h0e4e1: out <= 12'h603;
      20'h0e4e2: out <= 12'h603;
      20'h0e4e3: out <= 12'h603;
      20'h0e4e4: out <= 12'h603;
      20'h0e4e5: out <= 12'h603;
      20'h0e4e6: out <= 12'h603;
      20'h0e4e7: out <= 12'h603;
      20'h0e4e8: out <= 12'h603;
      20'h0e4e9: out <= 12'h603;
      20'h0e4ea: out <= 12'h603;
      20'h0e4eb: out <= 12'h603;
      20'h0e4ec: out <= 12'h603;
      20'h0e4ed: out <= 12'h603;
      20'h0e4ee: out <= 12'h603;
      20'h0e4ef: out <= 12'h603;
      20'h0e4f0: out <= 12'hfff;
      20'h0e4f1: out <= 12'hfff;
      20'h0e4f2: out <= 12'hc7f;
      20'h0e4f3: out <= 12'h000;
      20'h0e4f4: out <= 12'h000;
      20'h0e4f5: out <= 12'h000;
      20'h0e4f6: out <= 12'h000;
      20'h0e4f7: out <= 12'h000;
      20'h0e4f8: out <= 12'h000;
      20'h0e4f9: out <= 12'h000;
      20'h0e4fa: out <= 12'hc7f;
      20'h0e4fb: out <= 12'hc7f;
      20'h0e4fc: out <= 12'hc7f;
      20'h0e4fd: out <= 12'hc7f;
      20'h0e4fe: out <= 12'h000;
      20'h0e4ff: out <= 12'h000;
      20'h0e500: out <= 12'h000;
      20'h0e501: out <= 12'h000;
      20'h0e502: out <= 12'hc7f;
      20'h0e503: out <= 12'hc7f;
      20'h0e504: out <= 12'hc7f;
      20'h0e505: out <= 12'h000;
      20'h0e506: out <= 12'h000;
      20'h0e507: out <= 12'h000;
      20'h0e508: out <= 12'hc7f;
      20'h0e509: out <= 12'hc7f;
      20'h0e50a: out <= 12'hc7f;
      20'h0e50b: out <= 12'h000;
      20'h0e50c: out <= 12'h000;
      20'h0e50d: out <= 12'h000;
      20'h0e50e: out <= 12'hc7f;
      20'h0e50f: out <= 12'h000;
      20'h0e510: out <= 12'h000;
      20'h0e511: out <= 12'h000;
      20'h0e512: out <= 12'h000;
      20'h0e513: out <= 12'h000;
      20'h0e514: out <= 12'h000;
      20'h0e515: out <= 12'h000;
      20'h0e516: out <= 12'h72f;
      20'h0e517: out <= 12'h72f;
      20'h0e518: out <= 12'h603;
      20'h0e519: out <= 12'h603;
      20'h0e51a: out <= 12'h603;
      20'h0e51b: out <= 12'h603;
      20'h0e51c: out <= 12'h603;
      20'h0e51d: out <= 12'h603;
      20'h0e51e: out <= 12'h603;
      20'h0e51f: out <= 12'h603;
      20'h0e520: out <= 12'h603;
      20'h0e521: out <= 12'h603;
      20'h0e522: out <= 12'h603;
      20'h0e523: out <= 12'h603;
      20'h0e524: out <= 12'h603;
      20'h0e525: out <= 12'h603;
      20'h0e526: out <= 12'h603;
      20'h0e527: out <= 12'h603;
      20'h0e528: out <= 12'h603;
      20'h0e529: out <= 12'h603;
      20'h0e52a: out <= 12'h603;
      20'h0e52b: out <= 12'h603;
      20'h0e52c: out <= 12'h603;
      20'h0e52d: out <= 12'h603;
      20'h0e52e: out <= 12'h603;
      20'h0e52f: out <= 12'h603;
      20'h0e530: out <= 12'h603;
      20'h0e531: out <= 12'h603;
      20'h0e532: out <= 12'h603;
      20'h0e533: out <= 12'h603;
      20'h0e534: out <= 12'h603;
      20'h0e535: out <= 12'h603;
      20'h0e536: out <= 12'h603;
      20'h0e537: out <= 12'h603;
      20'h0e538: out <= 12'h603;
      20'h0e539: out <= 12'h603;
      20'h0e53a: out <= 12'h603;
      20'h0e53b: out <= 12'h603;
      20'h0e53c: out <= 12'h603;
      20'h0e53d: out <= 12'h603;
      20'h0e53e: out <= 12'h603;
      20'h0e53f: out <= 12'h603;
      20'h0e540: out <= 12'h603;
      20'h0e541: out <= 12'h603;
      20'h0e542: out <= 12'h603;
      20'h0e543: out <= 12'h603;
      20'h0e544: out <= 12'h603;
      20'h0e545: out <= 12'h603;
      20'h0e546: out <= 12'h603;
      20'h0e547: out <= 12'h603;
      20'h0e548: out <= 12'h603;
      20'h0e549: out <= 12'h603;
      20'h0e54a: out <= 12'h603;
      20'h0e54b: out <= 12'h603;
      20'h0e54c: out <= 12'h603;
      20'h0e54d: out <= 12'h603;
      20'h0e54e: out <= 12'h603;
      20'h0e54f: out <= 12'h603;
      20'h0e550: out <= 12'h603;
      20'h0e551: out <= 12'h603;
      20'h0e552: out <= 12'h603;
      20'h0e553: out <= 12'h603;
      20'h0e554: out <= 12'h603;
      20'h0e555: out <= 12'h603;
      20'h0e556: out <= 12'h603;
      20'h0e557: out <= 12'h603;
      20'h0e558: out <= 12'h603;
      20'h0e559: out <= 12'h603;
      20'h0e55a: out <= 12'h603;
      20'h0e55b: out <= 12'h603;
      20'h0e55c: out <= 12'h603;
      20'h0e55d: out <= 12'h603;
      20'h0e55e: out <= 12'h603;
      20'h0e55f: out <= 12'h603;
      20'h0e560: out <= 12'h603;
      20'h0e561: out <= 12'h603;
      20'h0e562: out <= 12'h603;
      20'h0e563: out <= 12'h603;
      20'h0e564: out <= 12'h603;
      20'h0e565: out <= 12'h603;
      20'h0e566: out <= 12'h603;
      20'h0e567: out <= 12'h603;
      20'h0e568: out <= 12'h603;
      20'h0e569: out <= 12'h603;
      20'h0e56a: out <= 12'h603;
      20'h0e56b: out <= 12'h603;
      20'h0e56c: out <= 12'h603;
      20'h0e56d: out <= 12'h603;
      20'h0e56e: out <= 12'h603;
      20'h0e56f: out <= 12'h603;
      20'h0e570: out <= 12'hee9;
      20'h0e571: out <= 12'hf87;
      20'h0e572: out <= 12'hf87;
      20'h0e573: out <= 12'hf87;
      20'h0e574: out <= 12'hf87;
      20'h0e575: out <= 12'hf87;
      20'h0e576: out <= 12'hf87;
      20'h0e577: out <= 12'hb27;
      20'h0e578: out <= 12'h000;
      20'h0e579: out <= 12'h000;
      20'h0e57a: out <= 12'h000;
      20'h0e57b: out <= 12'h000;
      20'h0e57c: out <= 12'h000;
      20'h0e57d: out <= 12'h000;
      20'h0e57e: out <= 12'h000;
      20'h0e57f: out <= 12'h000;
      20'h0e580: out <= 12'h000;
      20'h0e581: out <= 12'h000;
      20'h0e582: out <= 12'h000;
      20'h0e583: out <= 12'h666;
      20'h0e584: out <= 12'h666;
      20'h0e585: out <= 12'hfff;
      20'h0e586: out <= 12'h666;
      20'h0e587: out <= 12'hfff;
      20'h0e588: out <= 12'hbbb;
      20'h0e589: out <= 12'hbbb;
      20'h0e58a: out <= 12'h666;
      20'h0e58b: out <= 12'h666;
      20'h0e58c: out <= 12'h666;
      20'h0e58d: out <= 12'h666;
      20'h0e58e: out <= 12'h000;
      20'h0e58f: out <= 12'h000;
      20'h0e590: out <= 12'h000;
      20'h0e591: out <= 12'h000;
      20'h0e592: out <= 12'hbbb;
      20'h0e593: out <= 12'h000;
      20'h0e594: out <= 12'h000;
      20'h0e595: out <= 12'h000;
      20'h0e596: out <= 12'hbbb;
      20'h0e597: out <= 12'h000;
      20'h0e598: out <= 12'h999;
      20'h0e599: out <= 12'h999;
      20'h0e59a: out <= 12'h999;
      20'h0e59b: out <= 12'h999;
      20'h0e59c: out <= 12'h999;
      20'h0e59d: out <= 12'h999;
      20'h0e59e: out <= 12'h999;
      20'h0e59f: out <= 12'h999;
      20'h0e5a0: out <= 12'hbbb;
      20'h0e5a1: out <= 12'hbbb;
      20'h0e5a2: out <= 12'hbbb;
      20'h0e5a3: out <= 12'hbbb;
      20'h0e5a4: out <= 12'hbbb;
      20'h0e5a5: out <= 12'hbbb;
      20'h0e5a6: out <= 12'hbbb;
      20'h0e5a7: out <= 12'hbbb;
      20'h0e5a8: out <= 12'h000;
      20'h0e5a9: out <= 12'h000;
      20'h0e5aa: out <= 12'h000;
      20'h0e5ab: out <= 12'h000;
      20'h0e5ac: out <= 12'h000;
      20'h0e5ad: out <= 12'h000;
      20'h0e5ae: out <= 12'h000;
      20'h0e5af: out <= 12'h000;
      20'h0e5b0: out <= 12'hfff;
      20'h0e5b1: out <= 12'hfff;
      20'h0e5b2: out <= 12'hbbb;
      20'h0e5b3: out <= 12'hbbb;
      20'h0e5b4: out <= 12'hbbb;
      20'h0e5b5: out <= 12'hbbb;
      20'h0e5b6: out <= 12'hbbb;
      20'h0e5b7: out <= 12'hbbb;
      20'h0e5b8: out <= 12'hbbb;
      20'h0e5b9: out <= 12'hbbb;
      20'h0e5ba: out <= 12'hbbb;
      20'h0e5bb: out <= 12'hbbb;
      20'h0e5bc: out <= 12'hbbb;
      20'h0e5bd: out <= 12'hbbb;
      20'h0e5be: out <= 12'hbbb;
      20'h0e5bf: out <= 12'hbbb;
      20'h0e5c0: out <= 12'hbbb;
      20'h0e5c1: out <= 12'hbbb;
      20'h0e5c2: out <= 12'hbbb;
      20'h0e5c3: out <= 12'hbbb;
      20'h0e5c4: out <= 12'hbbb;
      20'h0e5c5: out <= 12'hbbb;
      20'h0e5c6: out <= 12'hbbb;
      20'h0e5c7: out <= 12'hbbb;
      20'h0e5c8: out <= 12'hbbb;
      20'h0e5c9: out <= 12'hbbb;
      20'h0e5ca: out <= 12'hbbb;
      20'h0e5cb: out <= 12'hbbb;
      20'h0e5cc: out <= 12'hbbb;
      20'h0e5cd: out <= 12'hbbb;
      20'h0e5ce: out <= 12'hbbb;
      20'h0e5cf: out <= 12'hbbb;
      20'h0e5d0: out <= 12'hbbb;
      20'h0e5d1: out <= 12'hbbb;
      20'h0e5d2: out <= 12'hbbb;
      20'h0e5d3: out <= 12'hbbb;
      20'h0e5d4: out <= 12'hbbb;
      20'h0e5d5: out <= 12'hbbb;
      20'h0e5d6: out <= 12'hbbb;
      20'h0e5d7: out <= 12'hbbb;
      20'h0e5d8: out <= 12'hbbb;
      20'h0e5d9: out <= 12'hbbb;
      20'h0e5da: out <= 12'hbbb;
      20'h0e5db: out <= 12'hbbb;
      20'h0e5dc: out <= 12'hbbb;
      20'h0e5dd: out <= 12'hbbb;
      20'h0e5de: out <= 12'h666;
      20'h0e5df: out <= 12'h666;
      20'h0e5e0: out <= 12'h603;
      20'h0e5e1: out <= 12'h603;
      20'h0e5e2: out <= 12'h603;
      20'h0e5e3: out <= 12'h603;
      20'h0e5e4: out <= 12'h603;
      20'h0e5e5: out <= 12'h603;
      20'h0e5e6: out <= 12'h603;
      20'h0e5e7: out <= 12'h603;
      20'h0e5e8: out <= 12'h603;
      20'h0e5e9: out <= 12'h603;
      20'h0e5ea: out <= 12'h603;
      20'h0e5eb: out <= 12'h603;
      20'h0e5ec: out <= 12'h603;
      20'h0e5ed: out <= 12'h603;
      20'h0e5ee: out <= 12'h603;
      20'h0e5ef: out <= 12'h603;
      20'h0e5f0: out <= 12'h603;
      20'h0e5f1: out <= 12'h603;
      20'h0e5f2: out <= 12'h603;
      20'h0e5f3: out <= 12'h603;
      20'h0e5f4: out <= 12'h603;
      20'h0e5f5: out <= 12'h603;
      20'h0e5f6: out <= 12'h603;
      20'h0e5f7: out <= 12'h603;
      20'h0e5f8: out <= 12'h603;
      20'h0e5f9: out <= 12'h603;
      20'h0e5fa: out <= 12'h603;
      20'h0e5fb: out <= 12'h603;
      20'h0e5fc: out <= 12'h603;
      20'h0e5fd: out <= 12'h603;
      20'h0e5fe: out <= 12'h603;
      20'h0e5ff: out <= 12'h603;
      20'h0e600: out <= 12'h603;
      20'h0e601: out <= 12'h603;
      20'h0e602: out <= 12'h603;
      20'h0e603: out <= 12'h603;
      20'h0e604: out <= 12'h603;
      20'h0e605: out <= 12'h603;
      20'h0e606: out <= 12'h603;
      20'h0e607: out <= 12'h603;
      20'h0e608: out <= 12'hfff;
      20'h0e609: out <= 12'hfff;
      20'h0e60a: out <= 12'h000;
      20'h0e60b: out <= 12'h000;
      20'h0e60c: out <= 12'h000;
      20'h0e60d: out <= 12'hc7f;
      20'h0e60e: out <= 12'hc7f;
      20'h0e60f: out <= 12'hc7f;
      20'h0e610: out <= 12'hc7f;
      20'h0e611: out <= 12'h000;
      20'h0e612: out <= 12'h000;
      20'h0e613: out <= 12'hc7f;
      20'h0e614: out <= 12'hc7f;
      20'h0e615: out <= 12'h000;
      20'h0e616: out <= 12'h000;
      20'h0e617: out <= 12'hc7f;
      20'h0e618: out <= 12'hc7f;
      20'h0e619: out <= 12'h000;
      20'h0e61a: out <= 12'h000;
      20'h0e61b: out <= 12'hc7f;
      20'h0e61c: out <= 12'hc7f;
      20'h0e61d: out <= 12'h000;
      20'h0e61e: out <= 12'h000;
      20'h0e61f: out <= 12'h000;
      20'h0e620: out <= 12'h000;
      20'h0e621: out <= 12'hc7f;
      20'h0e622: out <= 12'h000;
      20'h0e623: out <= 12'h000;
      20'h0e624: out <= 12'h000;
      20'h0e625: out <= 12'h000;
      20'h0e626: out <= 12'hc7f;
      20'h0e627: out <= 12'h000;
      20'h0e628: out <= 12'h000;
      20'h0e629: out <= 12'h000;
      20'h0e62a: out <= 12'hc7f;
      20'h0e62b: out <= 12'hc7f;
      20'h0e62c: out <= 12'hc7f;
      20'h0e62d: out <= 12'hc7f;
      20'h0e62e: out <= 12'h72f;
      20'h0e62f: out <= 12'h72f;
      20'h0e630: out <= 12'h603;
      20'h0e631: out <= 12'h603;
      20'h0e632: out <= 12'h603;
      20'h0e633: out <= 12'h603;
      20'h0e634: out <= 12'h603;
      20'h0e635: out <= 12'h603;
      20'h0e636: out <= 12'h603;
      20'h0e637: out <= 12'h603;
      20'h0e638: out <= 12'h603;
      20'h0e639: out <= 12'h603;
      20'h0e63a: out <= 12'h603;
      20'h0e63b: out <= 12'h603;
      20'h0e63c: out <= 12'h603;
      20'h0e63d: out <= 12'h603;
      20'h0e63e: out <= 12'h603;
      20'h0e63f: out <= 12'h603;
      20'h0e640: out <= 12'h603;
      20'h0e641: out <= 12'h603;
      20'h0e642: out <= 12'h603;
      20'h0e643: out <= 12'h603;
      20'h0e644: out <= 12'h603;
      20'h0e645: out <= 12'h603;
      20'h0e646: out <= 12'h603;
      20'h0e647: out <= 12'h603;
      20'h0e648: out <= 12'h603;
      20'h0e649: out <= 12'h603;
      20'h0e64a: out <= 12'h603;
      20'h0e64b: out <= 12'h603;
      20'h0e64c: out <= 12'h603;
      20'h0e64d: out <= 12'h603;
      20'h0e64e: out <= 12'h603;
      20'h0e64f: out <= 12'h603;
      20'h0e650: out <= 12'h603;
      20'h0e651: out <= 12'h603;
      20'h0e652: out <= 12'h603;
      20'h0e653: out <= 12'h603;
      20'h0e654: out <= 12'h603;
      20'h0e655: out <= 12'h603;
      20'h0e656: out <= 12'h603;
      20'h0e657: out <= 12'h603;
      20'h0e658: out <= 12'h603;
      20'h0e659: out <= 12'h603;
      20'h0e65a: out <= 12'h603;
      20'h0e65b: out <= 12'h603;
      20'h0e65c: out <= 12'h603;
      20'h0e65d: out <= 12'h603;
      20'h0e65e: out <= 12'h603;
      20'h0e65f: out <= 12'h603;
      20'h0e660: out <= 12'h603;
      20'h0e661: out <= 12'h603;
      20'h0e662: out <= 12'h603;
      20'h0e663: out <= 12'h603;
      20'h0e664: out <= 12'h603;
      20'h0e665: out <= 12'h603;
      20'h0e666: out <= 12'h603;
      20'h0e667: out <= 12'h603;
      20'h0e668: out <= 12'h603;
      20'h0e669: out <= 12'h603;
      20'h0e66a: out <= 12'h603;
      20'h0e66b: out <= 12'h603;
      20'h0e66c: out <= 12'h603;
      20'h0e66d: out <= 12'h603;
      20'h0e66e: out <= 12'h603;
      20'h0e66f: out <= 12'h603;
      20'h0e670: out <= 12'h603;
      20'h0e671: out <= 12'h603;
      20'h0e672: out <= 12'h603;
      20'h0e673: out <= 12'h603;
      20'h0e674: out <= 12'h603;
      20'h0e675: out <= 12'h603;
      20'h0e676: out <= 12'h603;
      20'h0e677: out <= 12'h603;
      20'h0e678: out <= 12'h603;
      20'h0e679: out <= 12'h603;
      20'h0e67a: out <= 12'h603;
      20'h0e67b: out <= 12'h603;
      20'h0e67c: out <= 12'h603;
      20'h0e67d: out <= 12'h603;
      20'h0e67e: out <= 12'h603;
      20'h0e67f: out <= 12'h603;
      20'h0e680: out <= 12'h603;
      20'h0e681: out <= 12'h603;
      20'h0e682: out <= 12'h603;
      20'h0e683: out <= 12'h603;
      20'h0e684: out <= 12'h603;
      20'h0e685: out <= 12'h603;
      20'h0e686: out <= 12'h603;
      20'h0e687: out <= 12'h603;
      20'h0e688: out <= 12'hee9;
      20'h0e689: out <= 12'hf87;
      20'h0e68a: out <= 12'hee9;
      20'h0e68b: out <= 12'hee9;
      20'h0e68c: out <= 12'hee9;
      20'h0e68d: out <= 12'hb27;
      20'h0e68e: out <= 12'hf87;
      20'h0e68f: out <= 12'hb27;
      20'h0e690: out <= 12'h000;
      20'h0e691: out <= 12'h000;
      20'h0e692: out <= 12'h000;
      20'h0e693: out <= 12'h000;
      20'h0e694: out <= 12'h000;
      20'h0e695: out <= 12'h000;
      20'h0e696: out <= 12'h000;
      20'h0e697: out <= 12'h000;
      20'h0e698: out <= 12'h000;
      20'h0e699: out <= 12'h000;
      20'h0e69a: out <= 12'h666;
      20'h0e69b: out <= 12'hbbb;
      20'h0e69c: out <= 12'h666;
      20'h0e69d: out <= 12'hfff;
      20'h0e69e: out <= 12'h666;
      20'h0e69f: out <= 12'hbbb;
      20'h0e6a0: out <= 12'hbbb;
      20'h0e6a1: out <= 12'h666;
      20'h0e6a2: out <= 12'h666;
      20'h0e6a3: out <= 12'h666;
      20'h0e6a4: out <= 12'h666;
      20'h0e6a5: out <= 12'hbbb;
      20'h0e6a6: out <= 12'h666;
      20'h0e6a7: out <= 12'h000;
      20'h0e6a8: out <= 12'h000;
      20'h0e6a9: out <= 12'h000;
      20'h0e6aa: out <= 12'h000;
      20'h0e6ab: out <= 12'hbbb;
      20'h0e6ac: out <= 12'h000;
      20'h0e6ad: out <= 12'hbbb;
      20'h0e6ae: out <= 12'h000;
      20'h0e6af: out <= 12'h000;
      20'h0e6b0: out <= 12'h999;
      20'h0e6b1: out <= 12'h999;
      20'h0e6b2: out <= 12'h999;
      20'h0e6b3: out <= 12'h999;
      20'h0e6b4: out <= 12'h999;
      20'h0e6b5: out <= 12'h999;
      20'h0e6b6: out <= 12'h999;
      20'h0e6b7: out <= 12'h999;
      20'h0e6b8: out <= 12'hbbb;
      20'h0e6b9: out <= 12'hbbb;
      20'h0e6ba: out <= 12'hbbb;
      20'h0e6bb: out <= 12'hbbb;
      20'h0e6bc: out <= 12'hbbb;
      20'h0e6bd: out <= 12'hbbb;
      20'h0e6be: out <= 12'hbbb;
      20'h0e6bf: out <= 12'hbbb;
      20'h0e6c0: out <= 12'h000;
      20'h0e6c1: out <= 12'h000;
      20'h0e6c2: out <= 12'h000;
      20'h0e6c3: out <= 12'h000;
      20'h0e6c4: out <= 12'h000;
      20'h0e6c5: out <= 12'h000;
      20'h0e6c6: out <= 12'h000;
      20'h0e6c7: out <= 12'h000;
      20'h0e6c8: out <= 12'hfff;
      20'h0e6c9: out <= 12'hfff;
      20'h0e6ca: out <= 12'hbbb;
      20'h0e6cb: out <= 12'h666;
      20'h0e6cc: out <= 12'h666;
      20'h0e6cd: out <= 12'h666;
      20'h0e6ce: out <= 12'h666;
      20'h0e6cf: out <= 12'h666;
      20'h0e6d0: out <= 12'h666;
      20'h0e6d1: out <= 12'h666;
      20'h0e6d2: out <= 12'hfff;
      20'h0e6d3: out <= 12'hfff;
      20'h0e6d4: out <= 12'hfff;
      20'h0e6d5: out <= 12'hfff;
      20'h0e6d6: out <= 12'h666;
      20'h0e6d7: out <= 12'h666;
      20'h0e6d8: out <= 12'h666;
      20'h0e6d9: out <= 12'h666;
      20'h0e6da: out <= 12'hfff;
      20'h0e6db: out <= 12'hfff;
      20'h0e6dc: out <= 12'hfff;
      20'h0e6dd: out <= 12'h666;
      20'h0e6de: out <= 12'h666;
      20'h0e6df: out <= 12'h666;
      20'h0e6e0: out <= 12'hfff;
      20'h0e6e1: out <= 12'h666;
      20'h0e6e2: out <= 12'h666;
      20'h0e6e3: out <= 12'h666;
      20'h0e6e4: out <= 12'hfff;
      20'h0e6e5: out <= 12'hfff;
      20'h0e6e6: out <= 12'hfff;
      20'h0e6e7: out <= 12'h666;
      20'h0e6e8: out <= 12'h666;
      20'h0e6e9: out <= 12'h666;
      20'h0e6ea: out <= 12'h666;
      20'h0e6eb: out <= 12'hfff;
      20'h0e6ec: out <= 12'hfff;
      20'h0e6ed: out <= 12'hfff;
      20'h0e6ee: out <= 12'h666;
      20'h0e6ef: out <= 12'h666;
      20'h0e6f0: out <= 12'h666;
      20'h0e6f1: out <= 12'h666;
      20'h0e6f2: out <= 12'h666;
      20'h0e6f3: out <= 12'h666;
      20'h0e6f4: out <= 12'h666;
      20'h0e6f5: out <= 12'hbbb;
      20'h0e6f6: out <= 12'h666;
      20'h0e6f7: out <= 12'h666;
      20'h0e6f8: out <= 12'h603;
      20'h0e6f9: out <= 12'h603;
      20'h0e6fa: out <= 12'h603;
      20'h0e6fb: out <= 12'h603;
      20'h0e6fc: out <= 12'h603;
      20'h0e6fd: out <= 12'h603;
      20'h0e6fe: out <= 12'h603;
      20'h0e6ff: out <= 12'h603;
      20'h0e700: out <= 12'h603;
      20'h0e701: out <= 12'h603;
      20'h0e702: out <= 12'h603;
      20'h0e703: out <= 12'h603;
      20'h0e704: out <= 12'h603;
      20'h0e705: out <= 12'h603;
      20'h0e706: out <= 12'h603;
      20'h0e707: out <= 12'h603;
      20'h0e708: out <= 12'h603;
      20'h0e709: out <= 12'h603;
      20'h0e70a: out <= 12'h603;
      20'h0e70b: out <= 12'h603;
      20'h0e70c: out <= 12'h603;
      20'h0e70d: out <= 12'h603;
      20'h0e70e: out <= 12'h603;
      20'h0e70f: out <= 12'h603;
      20'h0e710: out <= 12'h603;
      20'h0e711: out <= 12'h603;
      20'h0e712: out <= 12'h603;
      20'h0e713: out <= 12'h603;
      20'h0e714: out <= 12'h603;
      20'h0e715: out <= 12'h603;
      20'h0e716: out <= 12'h603;
      20'h0e717: out <= 12'h603;
      20'h0e718: out <= 12'h603;
      20'h0e719: out <= 12'h603;
      20'h0e71a: out <= 12'h603;
      20'h0e71b: out <= 12'h603;
      20'h0e71c: out <= 12'h603;
      20'h0e71d: out <= 12'h603;
      20'h0e71e: out <= 12'h603;
      20'h0e71f: out <= 12'h603;
      20'h0e720: out <= 12'hfff;
      20'h0e721: out <= 12'hfff;
      20'h0e722: out <= 12'h000;
      20'h0e723: out <= 12'h000;
      20'h0e724: out <= 12'h000;
      20'h0e725: out <= 12'hc7f;
      20'h0e726: out <= 12'hc7f;
      20'h0e727: out <= 12'hc7f;
      20'h0e728: out <= 12'hc7f;
      20'h0e729: out <= 12'hc7f;
      20'h0e72a: out <= 12'hc7f;
      20'h0e72b: out <= 12'hc7f;
      20'h0e72c: out <= 12'h000;
      20'h0e72d: out <= 12'h000;
      20'h0e72e: out <= 12'hc7f;
      20'h0e72f: out <= 12'hc7f;
      20'h0e730: out <= 12'hc7f;
      20'h0e731: out <= 12'hc7f;
      20'h0e732: out <= 12'h000;
      20'h0e733: out <= 12'h000;
      20'h0e734: out <= 12'hc7f;
      20'h0e735: out <= 12'h000;
      20'h0e736: out <= 12'h000;
      20'h0e737: out <= 12'h000;
      20'h0e738: out <= 12'h000;
      20'h0e739: out <= 12'h000;
      20'h0e73a: out <= 12'h000;
      20'h0e73b: out <= 12'h000;
      20'h0e73c: out <= 12'h000;
      20'h0e73d: out <= 12'h000;
      20'h0e73e: out <= 12'hc7f;
      20'h0e73f: out <= 12'h000;
      20'h0e740: out <= 12'h000;
      20'h0e741: out <= 12'h000;
      20'h0e742: out <= 12'h000;
      20'h0e743: out <= 12'h000;
      20'h0e744: out <= 12'hc7f;
      20'h0e745: out <= 12'hc7f;
      20'h0e746: out <= 12'h72f;
      20'h0e747: out <= 12'h72f;
      20'h0e748: out <= 12'h603;
      20'h0e749: out <= 12'h603;
      20'h0e74a: out <= 12'h603;
      20'h0e74b: out <= 12'h603;
      20'h0e74c: out <= 12'h603;
      20'h0e74d: out <= 12'h603;
      20'h0e74e: out <= 12'h603;
      20'h0e74f: out <= 12'h603;
      20'h0e750: out <= 12'h603;
      20'h0e751: out <= 12'h603;
      20'h0e752: out <= 12'h603;
      20'h0e753: out <= 12'h603;
      20'h0e754: out <= 12'h603;
      20'h0e755: out <= 12'h603;
      20'h0e756: out <= 12'h603;
      20'h0e757: out <= 12'h603;
      20'h0e758: out <= 12'h603;
      20'h0e759: out <= 12'h603;
      20'h0e75a: out <= 12'h603;
      20'h0e75b: out <= 12'h603;
      20'h0e75c: out <= 12'h603;
      20'h0e75d: out <= 12'h603;
      20'h0e75e: out <= 12'h603;
      20'h0e75f: out <= 12'h603;
      20'h0e760: out <= 12'h603;
      20'h0e761: out <= 12'h603;
      20'h0e762: out <= 12'h603;
      20'h0e763: out <= 12'h603;
      20'h0e764: out <= 12'h603;
      20'h0e765: out <= 12'h603;
      20'h0e766: out <= 12'h603;
      20'h0e767: out <= 12'h603;
      20'h0e768: out <= 12'h603;
      20'h0e769: out <= 12'h603;
      20'h0e76a: out <= 12'h603;
      20'h0e76b: out <= 12'h603;
      20'h0e76c: out <= 12'h603;
      20'h0e76d: out <= 12'h603;
      20'h0e76e: out <= 12'h603;
      20'h0e76f: out <= 12'h603;
      20'h0e770: out <= 12'h603;
      20'h0e771: out <= 12'h603;
      20'h0e772: out <= 12'h603;
      20'h0e773: out <= 12'h603;
      20'h0e774: out <= 12'h603;
      20'h0e775: out <= 12'h603;
      20'h0e776: out <= 12'h603;
      20'h0e777: out <= 12'h603;
      20'h0e778: out <= 12'h603;
      20'h0e779: out <= 12'h603;
      20'h0e77a: out <= 12'h603;
      20'h0e77b: out <= 12'h603;
      20'h0e77c: out <= 12'h603;
      20'h0e77d: out <= 12'h603;
      20'h0e77e: out <= 12'h603;
      20'h0e77f: out <= 12'h603;
      20'h0e780: out <= 12'h603;
      20'h0e781: out <= 12'h603;
      20'h0e782: out <= 12'h603;
      20'h0e783: out <= 12'h603;
      20'h0e784: out <= 12'h603;
      20'h0e785: out <= 12'h603;
      20'h0e786: out <= 12'h603;
      20'h0e787: out <= 12'h603;
      20'h0e788: out <= 12'h603;
      20'h0e789: out <= 12'h603;
      20'h0e78a: out <= 12'h603;
      20'h0e78b: out <= 12'h603;
      20'h0e78c: out <= 12'h603;
      20'h0e78d: out <= 12'h603;
      20'h0e78e: out <= 12'h603;
      20'h0e78f: out <= 12'h603;
      20'h0e790: out <= 12'h603;
      20'h0e791: out <= 12'h603;
      20'h0e792: out <= 12'h603;
      20'h0e793: out <= 12'h603;
      20'h0e794: out <= 12'h603;
      20'h0e795: out <= 12'h603;
      20'h0e796: out <= 12'h603;
      20'h0e797: out <= 12'h603;
      20'h0e798: out <= 12'h603;
      20'h0e799: out <= 12'h603;
      20'h0e79a: out <= 12'h603;
      20'h0e79b: out <= 12'h603;
      20'h0e79c: out <= 12'h603;
      20'h0e79d: out <= 12'h603;
      20'h0e79e: out <= 12'h603;
      20'h0e79f: out <= 12'h603;
      20'h0e7a0: out <= 12'hee9;
      20'h0e7a1: out <= 12'hf87;
      20'h0e7a2: out <= 12'hee9;
      20'h0e7a3: out <= 12'hf87;
      20'h0e7a4: out <= 12'hf87;
      20'h0e7a5: out <= 12'hb27;
      20'h0e7a6: out <= 12'hf87;
      20'h0e7a7: out <= 12'hb27;
      20'h0e7a8: out <= 12'h000;
      20'h0e7a9: out <= 12'h000;
      20'h0e7aa: out <= 12'h000;
      20'h0e7ab: out <= 12'h000;
      20'h0e7ac: out <= 12'h000;
      20'h0e7ad: out <= 12'h000;
      20'h0e7ae: out <= 12'h000;
      20'h0e7af: out <= 12'h000;
      20'h0e7b0: out <= 12'h000;
      20'h0e7b1: out <= 12'h000;
      20'h0e7b2: out <= 12'h000;
      20'h0e7b3: out <= 12'h666;
      20'h0e7b4: out <= 12'h666;
      20'h0e7b5: out <= 12'hfff;
      20'h0e7b6: out <= 12'hfff;
      20'h0e7b7: out <= 12'h666;
      20'h0e7b8: out <= 12'h666;
      20'h0e7b9: out <= 12'h666;
      20'h0e7ba: out <= 12'h666;
      20'h0e7bb: out <= 12'h666;
      20'h0e7bc: out <= 12'h666;
      20'h0e7bd: out <= 12'h666;
      20'h0e7be: out <= 12'h000;
      20'h0e7bf: out <= 12'h000;
      20'h0e7c0: out <= 12'h000;
      20'h0e7c1: out <= 12'h000;
      20'h0e7c2: out <= 12'h000;
      20'h0e7c3: out <= 12'h000;
      20'h0e7c4: out <= 12'hbbb;
      20'h0e7c5: out <= 12'h000;
      20'h0e7c6: out <= 12'h000;
      20'h0e7c7: out <= 12'h000;
      20'h0e7c8: out <= 12'h999;
      20'h0e7c9: out <= 12'h999;
      20'h0e7ca: out <= 12'h999;
      20'h0e7cb: out <= 12'h999;
      20'h0e7cc: out <= 12'h999;
      20'h0e7cd: out <= 12'h999;
      20'h0e7ce: out <= 12'h999;
      20'h0e7cf: out <= 12'h999;
      20'h0e7d0: out <= 12'hbbb;
      20'h0e7d1: out <= 12'hbbb;
      20'h0e7d2: out <= 12'hbbb;
      20'h0e7d3: out <= 12'hbbb;
      20'h0e7d4: out <= 12'hbbb;
      20'h0e7d5: out <= 12'hbbb;
      20'h0e7d6: out <= 12'hbbb;
      20'h0e7d7: out <= 12'hbbb;
      20'h0e7d8: out <= 12'h000;
      20'h0e7d9: out <= 12'h000;
      20'h0e7da: out <= 12'h000;
      20'h0e7db: out <= 12'h000;
      20'h0e7dc: out <= 12'h000;
      20'h0e7dd: out <= 12'h000;
      20'h0e7de: out <= 12'h000;
      20'h0e7df: out <= 12'h000;
      20'h0e7e0: out <= 12'hfff;
      20'h0e7e1: out <= 12'hfff;
      20'h0e7e2: out <= 12'hbbb;
      20'h0e7e3: out <= 12'h666;
      20'h0e7e4: out <= 12'h666;
      20'h0e7e5: out <= 12'h666;
      20'h0e7e6: out <= 12'h666;
      20'h0e7e7: out <= 12'h666;
      20'h0e7e8: out <= 12'h666;
      20'h0e7e9: out <= 12'h666;
      20'h0e7ea: out <= 12'h666;
      20'h0e7eb: out <= 12'hfff;
      20'h0e7ec: out <= 12'hfff;
      20'h0e7ed: out <= 12'h666;
      20'h0e7ee: out <= 12'h666;
      20'h0e7ef: out <= 12'h666;
      20'h0e7f0: out <= 12'h666;
      20'h0e7f1: out <= 12'h666;
      20'h0e7f2: out <= 12'h666;
      20'h0e7f3: out <= 12'hfff;
      20'h0e7f4: out <= 12'hfff;
      20'h0e7f5: out <= 12'h666;
      20'h0e7f6: out <= 12'h666;
      20'h0e7f7: out <= 12'h666;
      20'h0e7f8: out <= 12'hfff;
      20'h0e7f9: out <= 12'h666;
      20'h0e7fa: out <= 12'h666;
      20'h0e7fb: out <= 12'h666;
      20'h0e7fc: out <= 12'hfff;
      20'h0e7fd: out <= 12'hfff;
      20'h0e7fe: out <= 12'h666;
      20'h0e7ff: out <= 12'h666;
      20'h0e800: out <= 12'h666;
      20'h0e801: out <= 12'h666;
      20'h0e802: out <= 12'h666;
      20'h0e803: out <= 12'h666;
      20'h0e804: out <= 12'hfff;
      20'h0e805: out <= 12'hfff;
      20'h0e806: out <= 12'h666;
      20'h0e807: out <= 12'h666;
      20'h0e808: out <= 12'h666;
      20'h0e809: out <= 12'h666;
      20'h0e80a: out <= 12'h666;
      20'h0e80b: out <= 12'h666;
      20'h0e80c: out <= 12'h666;
      20'h0e80d: out <= 12'hbbb;
      20'h0e80e: out <= 12'h666;
      20'h0e80f: out <= 12'h666;
      20'h0e810: out <= 12'h603;
      20'h0e811: out <= 12'h603;
      20'h0e812: out <= 12'h603;
      20'h0e813: out <= 12'h603;
      20'h0e814: out <= 12'h603;
      20'h0e815: out <= 12'h603;
      20'h0e816: out <= 12'h603;
      20'h0e817: out <= 12'h603;
      20'h0e818: out <= 12'h603;
      20'h0e819: out <= 12'h603;
      20'h0e81a: out <= 12'h603;
      20'h0e81b: out <= 12'h603;
      20'h0e81c: out <= 12'h603;
      20'h0e81d: out <= 12'h603;
      20'h0e81e: out <= 12'h603;
      20'h0e81f: out <= 12'h603;
      20'h0e820: out <= 12'h603;
      20'h0e821: out <= 12'h603;
      20'h0e822: out <= 12'h603;
      20'h0e823: out <= 12'h603;
      20'h0e824: out <= 12'h603;
      20'h0e825: out <= 12'h603;
      20'h0e826: out <= 12'h603;
      20'h0e827: out <= 12'h603;
      20'h0e828: out <= 12'h603;
      20'h0e829: out <= 12'h603;
      20'h0e82a: out <= 12'h603;
      20'h0e82b: out <= 12'h603;
      20'h0e82c: out <= 12'h603;
      20'h0e82d: out <= 12'h603;
      20'h0e82e: out <= 12'h603;
      20'h0e82f: out <= 12'h603;
      20'h0e830: out <= 12'h603;
      20'h0e831: out <= 12'h603;
      20'h0e832: out <= 12'h603;
      20'h0e833: out <= 12'h603;
      20'h0e834: out <= 12'h603;
      20'h0e835: out <= 12'h603;
      20'h0e836: out <= 12'h603;
      20'h0e837: out <= 12'h603;
      20'h0e838: out <= 12'hfff;
      20'h0e839: out <= 12'hfff;
      20'h0e83a: out <= 12'h000;
      20'h0e83b: out <= 12'h000;
      20'h0e83c: out <= 12'h000;
      20'h0e83d: out <= 12'hc7f;
      20'h0e83e: out <= 12'hc7f;
      20'h0e83f: out <= 12'h000;
      20'h0e840: out <= 12'h000;
      20'h0e841: out <= 12'h000;
      20'h0e842: out <= 12'h000;
      20'h0e843: out <= 12'hc7f;
      20'h0e844: out <= 12'h000;
      20'h0e845: out <= 12'h000;
      20'h0e846: out <= 12'h000;
      20'h0e847: out <= 12'h000;
      20'h0e848: out <= 12'h000;
      20'h0e849: out <= 12'h000;
      20'h0e84a: out <= 12'h000;
      20'h0e84b: out <= 12'h000;
      20'h0e84c: out <= 12'hc7f;
      20'h0e84d: out <= 12'h000;
      20'h0e84e: out <= 12'h000;
      20'h0e84f: out <= 12'hc7f;
      20'h0e850: out <= 12'h000;
      20'h0e851: out <= 12'h000;
      20'h0e852: out <= 12'h000;
      20'h0e853: out <= 12'hc7f;
      20'h0e854: out <= 12'h000;
      20'h0e855: out <= 12'h000;
      20'h0e856: out <= 12'hc7f;
      20'h0e857: out <= 12'h000;
      20'h0e858: out <= 12'h000;
      20'h0e859: out <= 12'h000;
      20'h0e85a: out <= 12'hc7f;
      20'h0e85b: out <= 12'hc7f;
      20'h0e85c: out <= 12'hc7f;
      20'h0e85d: out <= 12'hc7f;
      20'h0e85e: out <= 12'h72f;
      20'h0e85f: out <= 12'h72f;
      20'h0e860: out <= 12'h603;
      20'h0e861: out <= 12'h603;
      20'h0e862: out <= 12'h603;
      20'h0e863: out <= 12'h603;
      20'h0e864: out <= 12'h603;
      20'h0e865: out <= 12'h603;
      20'h0e866: out <= 12'h603;
      20'h0e867: out <= 12'h603;
      20'h0e868: out <= 12'h603;
      20'h0e869: out <= 12'h603;
      20'h0e86a: out <= 12'h603;
      20'h0e86b: out <= 12'h603;
      20'h0e86c: out <= 12'h603;
      20'h0e86d: out <= 12'h603;
      20'h0e86e: out <= 12'h603;
      20'h0e86f: out <= 12'h603;
      20'h0e870: out <= 12'h603;
      20'h0e871: out <= 12'h603;
      20'h0e872: out <= 12'h603;
      20'h0e873: out <= 12'h603;
      20'h0e874: out <= 12'h603;
      20'h0e875: out <= 12'h603;
      20'h0e876: out <= 12'h603;
      20'h0e877: out <= 12'h603;
      20'h0e878: out <= 12'h603;
      20'h0e879: out <= 12'h603;
      20'h0e87a: out <= 12'h603;
      20'h0e87b: out <= 12'h603;
      20'h0e87c: out <= 12'h603;
      20'h0e87d: out <= 12'h603;
      20'h0e87e: out <= 12'h603;
      20'h0e87f: out <= 12'h603;
      20'h0e880: out <= 12'h603;
      20'h0e881: out <= 12'h603;
      20'h0e882: out <= 12'h603;
      20'h0e883: out <= 12'h603;
      20'h0e884: out <= 12'h603;
      20'h0e885: out <= 12'h603;
      20'h0e886: out <= 12'h603;
      20'h0e887: out <= 12'h603;
      20'h0e888: out <= 12'h603;
      20'h0e889: out <= 12'h603;
      20'h0e88a: out <= 12'h603;
      20'h0e88b: out <= 12'h603;
      20'h0e88c: out <= 12'h603;
      20'h0e88d: out <= 12'h603;
      20'h0e88e: out <= 12'h603;
      20'h0e88f: out <= 12'h603;
      20'h0e890: out <= 12'h603;
      20'h0e891: out <= 12'h603;
      20'h0e892: out <= 12'h603;
      20'h0e893: out <= 12'h603;
      20'h0e894: out <= 12'h603;
      20'h0e895: out <= 12'h603;
      20'h0e896: out <= 12'h603;
      20'h0e897: out <= 12'h603;
      20'h0e898: out <= 12'h603;
      20'h0e899: out <= 12'h603;
      20'h0e89a: out <= 12'h603;
      20'h0e89b: out <= 12'h603;
      20'h0e89c: out <= 12'h603;
      20'h0e89d: out <= 12'h603;
      20'h0e89e: out <= 12'h603;
      20'h0e89f: out <= 12'h603;
      20'h0e8a0: out <= 12'h603;
      20'h0e8a1: out <= 12'h603;
      20'h0e8a2: out <= 12'h603;
      20'h0e8a3: out <= 12'h603;
      20'h0e8a4: out <= 12'h603;
      20'h0e8a5: out <= 12'h603;
      20'h0e8a6: out <= 12'h603;
      20'h0e8a7: out <= 12'h603;
      20'h0e8a8: out <= 12'h603;
      20'h0e8a9: out <= 12'h603;
      20'h0e8aa: out <= 12'h603;
      20'h0e8ab: out <= 12'h603;
      20'h0e8ac: out <= 12'h603;
      20'h0e8ad: out <= 12'h603;
      20'h0e8ae: out <= 12'h603;
      20'h0e8af: out <= 12'h603;
      20'h0e8b0: out <= 12'h603;
      20'h0e8b1: out <= 12'h603;
      20'h0e8b2: out <= 12'h603;
      20'h0e8b3: out <= 12'h603;
      20'h0e8b4: out <= 12'h603;
      20'h0e8b5: out <= 12'h603;
      20'h0e8b6: out <= 12'h603;
      20'h0e8b7: out <= 12'h603;
      20'h0e8b8: out <= 12'hee9;
      20'h0e8b9: out <= 12'hf87;
      20'h0e8ba: out <= 12'hee9;
      20'h0e8bb: out <= 12'hf87;
      20'h0e8bc: out <= 12'hf87;
      20'h0e8bd: out <= 12'hb27;
      20'h0e8be: out <= 12'hf87;
      20'h0e8bf: out <= 12'hb27;
      20'h0e8c0: out <= 12'h000;
      20'h0e8c1: out <= 12'h000;
      20'h0e8c2: out <= 12'h000;
      20'h0e8c3: out <= 12'h000;
      20'h0e8c4: out <= 12'h000;
      20'h0e8c5: out <= 12'h000;
      20'h0e8c6: out <= 12'h000;
      20'h0e8c7: out <= 12'h000;
      20'h0e8c8: out <= 12'h000;
      20'h0e8c9: out <= 12'h000;
      20'h0e8ca: out <= 12'h666;
      20'h0e8cb: out <= 12'hbbb;
      20'h0e8cc: out <= 12'h666;
      20'h0e8cd: out <= 12'hfff;
      20'h0e8ce: out <= 12'hfff;
      20'h0e8cf: out <= 12'hbbb;
      20'h0e8d0: out <= 12'hbbb;
      20'h0e8d1: out <= 12'hbbb;
      20'h0e8d2: out <= 12'h666;
      20'h0e8d3: out <= 12'h666;
      20'h0e8d4: out <= 12'h666;
      20'h0e8d5: out <= 12'hbbb;
      20'h0e8d6: out <= 12'h666;
      20'h0e8d7: out <= 12'h000;
      20'h0e8d8: out <= 12'h000;
      20'h0e8d9: out <= 12'h000;
      20'h0e8da: out <= 12'h000;
      20'h0e8db: out <= 12'hbbb;
      20'h0e8dc: out <= 12'h000;
      20'h0e8dd: out <= 12'hbbb;
      20'h0e8de: out <= 12'h000;
      20'h0e8df: out <= 12'h000;
      20'h0e8e0: out <= 12'h999;
      20'h0e8e1: out <= 12'h999;
      20'h0e8e2: out <= 12'h999;
      20'h0e8e3: out <= 12'h999;
      20'h0e8e4: out <= 12'h999;
      20'h0e8e5: out <= 12'h999;
      20'h0e8e6: out <= 12'h999;
      20'h0e8e7: out <= 12'h999;
      20'h0e8e8: out <= 12'hbbb;
      20'h0e8e9: out <= 12'hbbb;
      20'h0e8ea: out <= 12'hbbb;
      20'h0e8eb: out <= 12'hbbb;
      20'h0e8ec: out <= 12'hbbb;
      20'h0e8ed: out <= 12'hbbb;
      20'h0e8ee: out <= 12'hbbb;
      20'h0e8ef: out <= 12'hbbb;
      20'h0e8f0: out <= 12'h000;
      20'h0e8f1: out <= 12'h000;
      20'h0e8f2: out <= 12'h000;
      20'h0e8f3: out <= 12'h000;
      20'h0e8f4: out <= 12'h000;
      20'h0e8f5: out <= 12'h000;
      20'h0e8f6: out <= 12'h000;
      20'h0e8f7: out <= 12'h000;
      20'h0e8f8: out <= 12'hfff;
      20'h0e8f9: out <= 12'hfff;
      20'h0e8fa: out <= 12'hbbb;
      20'h0e8fb: out <= 12'h666;
      20'h0e8fc: out <= 12'h666;
      20'h0e8fd: out <= 12'h666;
      20'h0e8fe: out <= 12'hfff;
      20'h0e8ff: out <= 12'hfff;
      20'h0e900: out <= 12'h666;
      20'h0e901: out <= 12'h666;
      20'h0e902: out <= 12'h666;
      20'h0e903: out <= 12'hfff;
      20'h0e904: out <= 12'h666;
      20'h0e905: out <= 12'h666;
      20'h0e906: out <= 12'h666;
      20'h0e907: out <= 12'hfff;
      20'h0e908: out <= 12'hfff;
      20'h0e909: out <= 12'h666;
      20'h0e90a: out <= 12'h666;
      20'h0e90b: out <= 12'h666;
      20'h0e90c: out <= 12'hfff;
      20'h0e90d: out <= 12'h666;
      20'h0e90e: out <= 12'h666;
      20'h0e90f: out <= 12'h666;
      20'h0e910: out <= 12'hfff;
      20'h0e911: out <= 12'h666;
      20'h0e912: out <= 12'h666;
      20'h0e913: out <= 12'h666;
      20'h0e914: out <= 12'hfff;
      20'h0e915: out <= 12'h666;
      20'h0e916: out <= 12'h666;
      20'h0e917: out <= 12'h666;
      20'h0e918: out <= 12'h666;
      20'h0e919: out <= 12'hfff;
      20'h0e91a: out <= 12'h666;
      20'h0e91b: out <= 12'h666;
      20'h0e91c: out <= 12'h666;
      20'h0e91d: out <= 12'hfff;
      20'h0e91e: out <= 12'h666;
      20'h0e91f: out <= 12'h666;
      20'h0e920: out <= 12'h666;
      20'h0e921: out <= 12'hfff;
      20'h0e922: out <= 12'hfff;
      20'h0e923: out <= 12'hfff;
      20'h0e924: out <= 12'hfff;
      20'h0e925: out <= 12'hbbb;
      20'h0e926: out <= 12'h666;
      20'h0e927: out <= 12'h666;
      20'h0e928: out <= 12'h603;
      20'h0e929: out <= 12'h603;
      20'h0e92a: out <= 12'h603;
      20'h0e92b: out <= 12'h603;
      20'h0e92c: out <= 12'h603;
      20'h0e92d: out <= 12'h603;
      20'h0e92e: out <= 12'h603;
      20'h0e92f: out <= 12'h603;
      20'h0e930: out <= 12'h603;
      20'h0e931: out <= 12'h603;
      20'h0e932: out <= 12'h603;
      20'h0e933: out <= 12'h603;
      20'h0e934: out <= 12'h603;
      20'h0e935: out <= 12'h603;
      20'h0e936: out <= 12'h603;
      20'h0e937: out <= 12'h603;
      20'h0e938: out <= 12'h603;
      20'h0e939: out <= 12'h603;
      20'h0e93a: out <= 12'h603;
      20'h0e93b: out <= 12'h603;
      20'h0e93c: out <= 12'h603;
      20'h0e93d: out <= 12'h603;
      20'h0e93e: out <= 12'h603;
      20'h0e93f: out <= 12'h603;
      20'h0e940: out <= 12'h603;
      20'h0e941: out <= 12'h603;
      20'h0e942: out <= 12'h603;
      20'h0e943: out <= 12'h603;
      20'h0e944: out <= 12'h603;
      20'h0e945: out <= 12'h603;
      20'h0e946: out <= 12'h603;
      20'h0e947: out <= 12'h603;
      20'h0e948: out <= 12'h603;
      20'h0e949: out <= 12'h603;
      20'h0e94a: out <= 12'h603;
      20'h0e94b: out <= 12'h603;
      20'h0e94c: out <= 12'h603;
      20'h0e94d: out <= 12'h603;
      20'h0e94e: out <= 12'h603;
      20'h0e94f: out <= 12'h603;
      20'h0e950: out <= 12'hfff;
      20'h0e951: out <= 12'hfff;
      20'h0e952: out <= 12'h000;
      20'h0e953: out <= 12'h000;
      20'h0e954: out <= 12'h000;
      20'h0e955: out <= 12'hc7f;
      20'h0e956: out <= 12'hc7f;
      20'h0e957: out <= 12'hc7f;
      20'h0e958: out <= 12'hc7f;
      20'h0e959: out <= 12'h000;
      20'h0e95a: out <= 12'h000;
      20'h0e95b: out <= 12'hc7f;
      20'h0e95c: out <= 12'h000;
      20'h0e95d: out <= 12'h000;
      20'h0e95e: out <= 12'hc7f;
      20'h0e95f: out <= 12'hc7f;
      20'h0e960: out <= 12'hc7f;
      20'h0e961: out <= 12'hc7f;
      20'h0e962: out <= 12'h000;
      20'h0e963: out <= 12'h000;
      20'h0e964: out <= 12'hc7f;
      20'h0e965: out <= 12'h000;
      20'h0e966: out <= 12'h000;
      20'h0e967: out <= 12'hc7f;
      20'h0e968: out <= 12'hc7f;
      20'h0e969: out <= 12'h000;
      20'h0e96a: out <= 12'hc7f;
      20'h0e96b: out <= 12'hc7f;
      20'h0e96c: out <= 12'h000;
      20'h0e96d: out <= 12'h000;
      20'h0e96e: out <= 12'hc7f;
      20'h0e96f: out <= 12'h000;
      20'h0e970: out <= 12'h000;
      20'h0e971: out <= 12'h000;
      20'h0e972: out <= 12'hc7f;
      20'h0e973: out <= 12'hc7f;
      20'h0e974: out <= 12'hc7f;
      20'h0e975: out <= 12'hc7f;
      20'h0e976: out <= 12'h72f;
      20'h0e977: out <= 12'h72f;
      20'h0e978: out <= 12'h603;
      20'h0e979: out <= 12'h603;
      20'h0e97a: out <= 12'h603;
      20'h0e97b: out <= 12'h603;
      20'h0e97c: out <= 12'h603;
      20'h0e97d: out <= 12'h603;
      20'h0e97e: out <= 12'h603;
      20'h0e97f: out <= 12'h603;
      20'h0e980: out <= 12'h603;
      20'h0e981: out <= 12'h603;
      20'h0e982: out <= 12'h603;
      20'h0e983: out <= 12'h603;
      20'h0e984: out <= 12'h603;
      20'h0e985: out <= 12'h603;
      20'h0e986: out <= 12'h603;
      20'h0e987: out <= 12'h603;
      20'h0e988: out <= 12'h603;
      20'h0e989: out <= 12'h603;
      20'h0e98a: out <= 12'h603;
      20'h0e98b: out <= 12'h603;
      20'h0e98c: out <= 12'h603;
      20'h0e98d: out <= 12'h603;
      20'h0e98e: out <= 12'h603;
      20'h0e98f: out <= 12'h603;
      20'h0e990: out <= 12'h603;
      20'h0e991: out <= 12'h603;
      20'h0e992: out <= 12'h603;
      20'h0e993: out <= 12'h603;
      20'h0e994: out <= 12'h603;
      20'h0e995: out <= 12'h603;
      20'h0e996: out <= 12'h603;
      20'h0e997: out <= 12'h603;
      20'h0e998: out <= 12'h603;
      20'h0e999: out <= 12'h603;
      20'h0e99a: out <= 12'h603;
      20'h0e99b: out <= 12'h603;
      20'h0e99c: out <= 12'h603;
      20'h0e99d: out <= 12'h603;
      20'h0e99e: out <= 12'h603;
      20'h0e99f: out <= 12'h603;
      20'h0e9a0: out <= 12'h603;
      20'h0e9a1: out <= 12'h603;
      20'h0e9a2: out <= 12'h603;
      20'h0e9a3: out <= 12'h603;
      20'h0e9a4: out <= 12'h603;
      20'h0e9a5: out <= 12'h603;
      20'h0e9a6: out <= 12'h603;
      20'h0e9a7: out <= 12'h603;
      20'h0e9a8: out <= 12'h603;
      20'h0e9a9: out <= 12'h603;
      20'h0e9aa: out <= 12'h603;
      20'h0e9ab: out <= 12'h603;
      20'h0e9ac: out <= 12'h603;
      20'h0e9ad: out <= 12'h603;
      20'h0e9ae: out <= 12'h603;
      20'h0e9af: out <= 12'h603;
      20'h0e9b0: out <= 12'h603;
      20'h0e9b1: out <= 12'h603;
      20'h0e9b2: out <= 12'h603;
      20'h0e9b3: out <= 12'h603;
      20'h0e9b4: out <= 12'h603;
      20'h0e9b5: out <= 12'h603;
      20'h0e9b6: out <= 12'h603;
      20'h0e9b7: out <= 12'h603;
      20'h0e9b8: out <= 12'h603;
      20'h0e9b9: out <= 12'h603;
      20'h0e9ba: out <= 12'h603;
      20'h0e9bb: out <= 12'h603;
      20'h0e9bc: out <= 12'h603;
      20'h0e9bd: out <= 12'h603;
      20'h0e9be: out <= 12'h603;
      20'h0e9bf: out <= 12'h603;
      20'h0e9c0: out <= 12'h603;
      20'h0e9c1: out <= 12'h603;
      20'h0e9c2: out <= 12'h603;
      20'h0e9c3: out <= 12'h603;
      20'h0e9c4: out <= 12'h603;
      20'h0e9c5: out <= 12'h603;
      20'h0e9c6: out <= 12'h603;
      20'h0e9c7: out <= 12'h603;
      20'h0e9c8: out <= 12'h603;
      20'h0e9c9: out <= 12'h603;
      20'h0e9ca: out <= 12'h603;
      20'h0e9cb: out <= 12'h603;
      20'h0e9cc: out <= 12'h603;
      20'h0e9cd: out <= 12'h603;
      20'h0e9ce: out <= 12'h603;
      20'h0e9cf: out <= 12'h603;
      20'h0e9d0: out <= 12'hee9;
      20'h0e9d1: out <= 12'hf87;
      20'h0e9d2: out <= 12'hee9;
      20'h0e9d3: out <= 12'hb27;
      20'h0e9d4: out <= 12'hb27;
      20'h0e9d5: out <= 12'hb27;
      20'h0e9d6: out <= 12'hf87;
      20'h0e9d7: out <= 12'hb27;
      20'h0e9d8: out <= 12'h000;
      20'h0e9d9: out <= 12'h000;
      20'h0e9da: out <= 12'h000;
      20'h0e9db: out <= 12'h000;
      20'h0e9dc: out <= 12'h000;
      20'h0e9dd: out <= 12'h000;
      20'h0e9de: out <= 12'h000;
      20'h0e9df: out <= 12'h000;
      20'h0e9e0: out <= 12'h000;
      20'h0e9e1: out <= 12'h000;
      20'h0e9e2: out <= 12'h000;
      20'h0e9e3: out <= 12'hbbb;
      20'h0e9e4: out <= 12'h000;
      20'h0e9e5: out <= 12'h666;
      20'h0e9e6: out <= 12'hfff;
      20'h0e9e7: out <= 12'hbbb;
      20'h0e9e8: out <= 12'hbbb;
      20'h0e9e9: out <= 12'hbbb;
      20'h0e9ea: out <= 12'h666;
      20'h0e9eb: out <= 12'h666;
      20'h0e9ec: out <= 12'h000;
      20'h0e9ed: out <= 12'hbbb;
      20'h0e9ee: out <= 12'h000;
      20'h0e9ef: out <= 12'h000;
      20'h0e9f0: out <= 12'h000;
      20'h0e9f1: out <= 12'h000;
      20'h0e9f2: out <= 12'hbbb;
      20'h0e9f3: out <= 12'h000;
      20'h0e9f4: out <= 12'h000;
      20'h0e9f5: out <= 12'h000;
      20'h0e9f6: out <= 12'hbbb;
      20'h0e9f7: out <= 12'h000;
      20'h0e9f8: out <= 12'h999;
      20'h0e9f9: out <= 12'h999;
      20'h0e9fa: out <= 12'h999;
      20'h0e9fb: out <= 12'h999;
      20'h0e9fc: out <= 12'h999;
      20'h0e9fd: out <= 12'h999;
      20'h0e9fe: out <= 12'h999;
      20'h0e9ff: out <= 12'h999;
      20'h0ea00: out <= 12'hbbb;
      20'h0ea01: out <= 12'hbbb;
      20'h0ea02: out <= 12'hbbb;
      20'h0ea03: out <= 12'hbbb;
      20'h0ea04: out <= 12'hbbb;
      20'h0ea05: out <= 12'hbbb;
      20'h0ea06: out <= 12'hbbb;
      20'h0ea07: out <= 12'hbbb;
      20'h0ea08: out <= 12'h000;
      20'h0ea09: out <= 12'h000;
      20'h0ea0a: out <= 12'h000;
      20'h0ea0b: out <= 12'h000;
      20'h0ea0c: out <= 12'h000;
      20'h0ea0d: out <= 12'h000;
      20'h0ea0e: out <= 12'h000;
      20'h0ea0f: out <= 12'h000;
      20'h0ea10: out <= 12'hfff;
      20'h0ea11: out <= 12'hfff;
      20'h0ea12: out <= 12'hbbb;
      20'h0ea13: out <= 12'h666;
      20'h0ea14: out <= 12'h666;
      20'h0ea15: out <= 12'h666;
      20'h0ea16: out <= 12'hfff;
      20'h0ea17: out <= 12'hfff;
      20'h0ea18: out <= 12'h666;
      20'h0ea19: out <= 12'h666;
      20'h0ea1a: out <= 12'h666;
      20'h0ea1b: out <= 12'hfff;
      20'h0ea1c: out <= 12'h666;
      20'h0ea1d: out <= 12'h666;
      20'h0ea1e: out <= 12'h666;
      20'h0ea1f: out <= 12'hfff;
      20'h0ea20: out <= 12'hfff;
      20'h0ea21: out <= 12'h666;
      20'h0ea22: out <= 12'h666;
      20'h0ea23: out <= 12'h666;
      20'h0ea24: out <= 12'hfff;
      20'h0ea25: out <= 12'h666;
      20'h0ea26: out <= 12'h666;
      20'h0ea27: out <= 12'h666;
      20'h0ea28: out <= 12'hfff;
      20'h0ea29: out <= 12'h666;
      20'h0ea2a: out <= 12'h666;
      20'h0ea2b: out <= 12'h666;
      20'h0ea2c: out <= 12'hfff;
      20'h0ea2d: out <= 12'h666;
      20'h0ea2e: out <= 12'h666;
      20'h0ea2f: out <= 12'h666;
      20'h0ea30: out <= 12'h666;
      20'h0ea31: out <= 12'hfff;
      20'h0ea32: out <= 12'hfff;
      20'h0ea33: out <= 12'hfff;
      20'h0ea34: out <= 12'hfff;
      20'h0ea35: out <= 12'hfff;
      20'h0ea36: out <= 12'h666;
      20'h0ea37: out <= 12'h666;
      20'h0ea38: out <= 12'h666;
      20'h0ea39: out <= 12'hfff;
      20'h0ea3a: out <= 12'hfff;
      20'h0ea3b: out <= 12'hfff;
      20'h0ea3c: out <= 12'hfff;
      20'h0ea3d: out <= 12'hbbb;
      20'h0ea3e: out <= 12'h666;
      20'h0ea3f: out <= 12'h666;
      20'h0ea40: out <= 12'h603;
      20'h0ea41: out <= 12'h603;
      20'h0ea42: out <= 12'h603;
      20'h0ea43: out <= 12'h603;
      20'h0ea44: out <= 12'h603;
      20'h0ea45: out <= 12'h603;
      20'h0ea46: out <= 12'h603;
      20'h0ea47: out <= 12'h603;
      20'h0ea48: out <= 12'h603;
      20'h0ea49: out <= 12'h603;
      20'h0ea4a: out <= 12'h603;
      20'h0ea4b: out <= 12'h603;
      20'h0ea4c: out <= 12'h603;
      20'h0ea4d: out <= 12'h603;
      20'h0ea4e: out <= 12'h603;
      20'h0ea4f: out <= 12'h603;
      20'h0ea50: out <= 12'h603;
      20'h0ea51: out <= 12'h603;
      20'h0ea52: out <= 12'h603;
      20'h0ea53: out <= 12'h603;
      20'h0ea54: out <= 12'h603;
      20'h0ea55: out <= 12'h603;
      20'h0ea56: out <= 12'h603;
      20'h0ea57: out <= 12'h603;
      20'h0ea58: out <= 12'h603;
      20'h0ea59: out <= 12'h603;
      20'h0ea5a: out <= 12'h603;
      20'h0ea5b: out <= 12'h603;
      20'h0ea5c: out <= 12'h603;
      20'h0ea5d: out <= 12'h603;
      20'h0ea5e: out <= 12'h603;
      20'h0ea5f: out <= 12'h603;
      20'h0ea60: out <= 12'h603;
      20'h0ea61: out <= 12'h603;
      20'h0ea62: out <= 12'h603;
      20'h0ea63: out <= 12'h603;
      20'h0ea64: out <= 12'h603;
      20'h0ea65: out <= 12'h603;
      20'h0ea66: out <= 12'h603;
      20'h0ea67: out <= 12'h603;
      20'h0ea68: out <= 12'hfff;
      20'h0ea69: out <= 12'hfff;
      20'h0ea6a: out <= 12'hc7f;
      20'h0ea6b: out <= 12'h000;
      20'h0ea6c: out <= 12'h000;
      20'h0ea6d: out <= 12'h000;
      20'h0ea6e: out <= 12'h000;
      20'h0ea6f: out <= 12'h000;
      20'h0ea70: out <= 12'h000;
      20'h0ea71: out <= 12'h000;
      20'h0ea72: out <= 12'hc7f;
      20'h0ea73: out <= 12'hc7f;
      20'h0ea74: out <= 12'h000;
      20'h0ea75: out <= 12'h000;
      20'h0ea76: out <= 12'hc7f;
      20'h0ea77: out <= 12'hc7f;
      20'h0ea78: out <= 12'hc7f;
      20'h0ea79: out <= 12'hc7f;
      20'h0ea7a: out <= 12'h000;
      20'h0ea7b: out <= 12'h000;
      20'h0ea7c: out <= 12'hc7f;
      20'h0ea7d: out <= 12'h000;
      20'h0ea7e: out <= 12'h000;
      20'h0ea7f: out <= 12'hc7f;
      20'h0ea80: out <= 12'hc7f;
      20'h0ea81: out <= 12'hc7f;
      20'h0ea82: out <= 12'hc7f;
      20'h0ea83: out <= 12'hc7f;
      20'h0ea84: out <= 12'h000;
      20'h0ea85: out <= 12'h000;
      20'h0ea86: out <= 12'hc7f;
      20'h0ea87: out <= 12'h000;
      20'h0ea88: out <= 12'h000;
      20'h0ea89: out <= 12'h000;
      20'h0ea8a: out <= 12'h000;
      20'h0ea8b: out <= 12'h000;
      20'h0ea8c: out <= 12'h000;
      20'h0ea8d: out <= 12'h000;
      20'h0ea8e: out <= 12'h72f;
      20'h0ea8f: out <= 12'h72f;
      20'h0ea90: out <= 12'h603;
      20'h0ea91: out <= 12'h603;
      20'h0ea92: out <= 12'h603;
      20'h0ea93: out <= 12'h603;
      20'h0ea94: out <= 12'h603;
      20'h0ea95: out <= 12'h603;
      20'h0ea96: out <= 12'h603;
      20'h0ea97: out <= 12'h603;
      20'h0ea98: out <= 12'h603;
      20'h0ea99: out <= 12'h603;
      20'h0ea9a: out <= 12'h603;
      20'h0ea9b: out <= 12'h603;
      20'h0ea9c: out <= 12'h603;
      20'h0ea9d: out <= 12'h603;
      20'h0ea9e: out <= 12'h603;
      20'h0ea9f: out <= 12'h603;
      20'h0eaa0: out <= 12'h603;
      20'h0eaa1: out <= 12'h603;
      20'h0eaa2: out <= 12'h603;
      20'h0eaa3: out <= 12'h603;
      20'h0eaa4: out <= 12'h603;
      20'h0eaa5: out <= 12'h603;
      20'h0eaa6: out <= 12'h603;
      20'h0eaa7: out <= 12'h603;
      20'h0eaa8: out <= 12'h603;
      20'h0eaa9: out <= 12'h603;
      20'h0eaaa: out <= 12'h603;
      20'h0eaab: out <= 12'h603;
      20'h0eaac: out <= 12'h603;
      20'h0eaad: out <= 12'h603;
      20'h0eaae: out <= 12'h603;
      20'h0eaaf: out <= 12'h603;
      20'h0eab0: out <= 12'h603;
      20'h0eab1: out <= 12'h603;
      20'h0eab2: out <= 12'h603;
      20'h0eab3: out <= 12'h603;
      20'h0eab4: out <= 12'h603;
      20'h0eab5: out <= 12'h603;
      20'h0eab6: out <= 12'h603;
      20'h0eab7: out <= 12'h603;
      20'h0eab8: out <= 12'h603;
      20'h0eab9: out <= 12'h603;
      20'h0eaba: out <= 12'h603;
      20'h0eabb: out <= 12'h603;
      20'h0eabc: out <= 12'h603;
      20'h0eabd: out <= 12'h603;
      20'h0eabe: out <= 12'h603;
      20'h0eabf: out <= 12'h603;
      20'h0eac0: out <= 12'h603;
      20'h0eac1: out <= 12'h603;
      20'h0eac2: out <= 12'h603;
      20'h0eac3: out <= 12'h603;
      20'h0eac4: out <= 12'h603;
      20'h0eac5: out <= 12'h603;
      20'h0eac6: out <= 12'h603;
      20'h0eac7: out <= 12'h603;
      20'h0eac8: out <= 12'h603;
      20'h0eac9: out <= 12'h603;
      20'h0eaca: out <= 12'h603;
      20'h0eacb: out <= 12'h603;
      20'h0eacc: out <= 12'h603;
      20'h0eacd: out <= 12'h603;
      20'h0eace: out <= 12'h603;
      20'h0eacf: out <= 12'h603;
      20'h0ead0: out <= 12'h603;
      20'h0ead1: out <= 12'h603;
      20'h0ead2: out <= 12'h603;
      20'h0ead3: out <= 12'h603;
      20'h0ead4: out <= 12'h603;
      20'h0ead5: out <= 12'h603;
      20'h0ead6: out <= 12'h603;
      20'h0ead7: out <= 12'h603;
      20'h0ead8: out <= 12'h603;
      20'h0ead9: out <= 12'h603;
      20'h0eada: out <= 12'h603;
      20'h0eadb: out <= 12'h603;
      20'h0eadc: out <= 12'h603;
      20'h0eadd: out <= 12'h603;
      20'h0eade: out <= 12'h603;
      20'h0eadf: out <= 12'h603;
      20'h0eae0: out <= 12'h603;
      20'h0eae1: out <= 12'h603;
      20'h0eae2: out <= 12'h603;
      20'h0eae3: out <= 12'h603;
      20'h0eae4: out <= 12'h603;
      20'h0eae5: out <= 12'h603;
      20'h0eae6: out <= 12'h603;
      20'h0eae7: out <= 12'h603;
      20'h0eae8: out <= 12'hee9;
      20'h0eae9: out <= 12'hf87;
      20'h0eaea: out <= 12'hf87;
      20'h0eaeb: out <= 12'hf87;
      20'h0eaec: out <= 12'hf87;
      20'h0eaed: out <= 12'hf87;
      20'h0eaee: out <= 12'hf87;
      20'h0eaef: out <= 12'hb27;
      20'h0eaf0: out <= 12'h000;
      20'h0eaf1: out <= 12'h000;
      20'h0eaf2: out <= 12'h000;
      20'h0eaf3: out <= 12'h000;
      20'h0eaf4: out <= 12'h000;
      20'h0eaf5: out <= 12'h000;
      20'h0eaf6: out <= 12'h000;
      20'h0eaf7: out <= 12'h000;
      20'h0eaf8: out <= 12'h000;
      20'h0eaf9: out <= 12'h000;
      20'h0eafa: out <= 12'h000;
      20'h0eafb: out <= 12'h000;
      20'h0eafc: out <= 12'h000;
      20'h0eafd: out <= 12'h000;
      20'h0eafe: out <= 12'h666;
      20'h0eaff: out <= 12'h666;
      20'h0eb00: out <= 12'h666;
      20'h0eb01: out <= 12'h666;
      20'h0eb02: out <= 12'h666;
      20'h0eb03: out <= 12'h000;
      20'h0eb04: out <= 12'h000;
      20'h0eb05: out <= 12'h000;
      20'h0eb06: out <= 12'h000;
      20'h0eb07: out <= 12'h000;
      20'h0eb08: out <= 12'h000;
      20'h0eb09: out <= 12'h000;
      20'h0eb0a: out <= 12'h000;
      20'h0eb0b: out <= 12'h000;
      20'h0eb0c: out <= 12'h000;
      20'h0eb0d: out <= 12'h000;
      20'h0eb0e: out <= 12'h000;
      20'h0eb0f: out <= 12'h000;
      20'h0eb10: out <= 12'h999;
      20'h0eb11: out <= 12'h999;
      20'h0eb12: out <= 12'h999;
      20'h0eb13: out <= 12'h999;
      20'h0eb14: out <= 12'h999;
      20'h0eb15: out <= 12'h999;
      20'h0eb16: out <= 12'h999;
      20'h0eb17: out <= 12'h999;
      20'h0eb18: out <= 12'hbbb;
      20'h0eb19: out <= 12'hbbb;
      20'h0eb1a: out <= 12'hbbb;
      20'h0eb1b: out <= 12'hbbb;
      20'h0eb1c: out <= 12'hbbb;
      20'h0eb1d: out <= 12'hbbb;
      20'h0eb1e: out <= 12'hbbb;
      20'h0eb1f: out <= 12'hbbb;
      20'h0eb20: out <= 12'h000;
      20'h0eb21: out <= 12'h000;
      20'h0eb22: out <= 12'h000;
      20'h0eb23: out <= 12'h000;
      20'h0eb24: out <= 12'h000;
      20'h0eb25: out <= 12'h000;
      20'h0eb26: out <= 12'h000;
      20'h0eb27: out <= 12'h000;
      20'h0eb28: out <= 12'hfff;
      20'h0eb29: out <= 12'hfff;
      20'h0eb2a: out <= 12'hbbb;
      20'h0eb2b: out <= 12'h666;
      20'h0eb2c: out <= 12'h666;
      20'h0eb2d: out <= 12'h666;
      20'h0eb2e: out <= 12'hfff;
      20'h0eb2f: out <= 12'hfff;
      20'h0eb30: out <= 12'h666;
      20'h0eb31: out <= 12'h666;
      20'h0eb32: out <= 12'h666;
      20'h0eb33: out <= 12'hfff;
      20'h0eb34: out <= 12'h666;
      20'h0eb35: out <= 12'h666;
      20'h0eb36: out <= 12'h666;
      20'h0eb37: out <= 12'hfff;
      20'h0eb38: out <= 12'hfff;
      20'h0eb39: out <= 12'h666;
      20'h0eb3a: out <= 12'h666;
      20'h0eb3b: out <= 12'h666;
      20'h0eb3c: out <= 12'hfff;
      20'h0eb3d: out <= 12'h666;
      20'h0eb3e: out <= 12'h666;
      20'h0eb3f: out <= 12'h666;
      20'h0eb40: out <= 12'hfff;
      20'h0eb41: out <= 12'h666;
      20'h0eb42: out <= 12'h666;
      20'h0eb43: out <= 12'h666;
      20'h0eb44: out <= 12'hfff;
      20'h0eb45: out <= 12'hfff;
      20'h0eb46: out <= 12'h666;
      20'h0eb47: out <= 12'h666;
      20'h0eb48: out <= 12'h666;
      20'h0eb49: out <= 12'h666;
      20'h0eb4a: out <= 12'h666;
      20'h0eb4b: out <= 12'hfff;
      20'h0eb4c: out <= 12'hfff;
      20'h0eb4d: out <= 12'hfff;
      20'h0eb4e: out <= 12'h666;
      20'h0eb4f: out <= 12'h666;
      20'h0eb50: out <= 12'h666;
      20'h0eb51: out <= 12'h666;
      20'h0eb52: out <= 12'h666;
      20'h0eb53: out <= 12'h666;
      20'h0eb54: out <= 12'hfff;
      20'h0eb55: out <= 12'hbbb;
      20'h0eb56: out <= 12'h666;
      20'h0eb57: out <= 12'h666;
      20'h0eb58: out <= 12'h603;
      20'h0eb59: out <= 12'h603;
      20'h0eb5a: out <= 12'h603;
      20'h0eb5b: out <= 12'h603;
      20'h0eb5c: out <= 12'h603;
      20'h0eb5d: out <= 12'h603;
      20'h0eb5e: out <= 12'h603;
      20'h0eb5f: out <= 12'h603;
      20'h0eb60: out <= 12'h603;
      20'h0eb61: out <= 12'h603;
      20'h0eb62: out <= 12'h603;
      20'h0eb63: out <= 12'h603;
      20'h0eb64: out <= 12'h603;
      20'h0eb65: out <= 12'h603;
      20'h0eb66: out <= 12'h603;
      20'h0eb67: out <= 12'h603;
      20'h0eb68: out <= 12'h603;
      20'h0eb69: out <= 12'h603;
      20'h0eb6a: out <= 12'h603;
      20'h0eb6b: out <= 12'h603;
      20'h0eb6c: out <= 12'h603;
      20'h0eb6d: out <= 12'h603;
      20'h0eb6e: out <= 12'h603;
      20'h0eb6f: out <= 12'h603;
      20'h0eb70: out <= 12'h603;
      20'h0eb71: out <= 12'h603;
      20'h0eb72: out <= 12'h603;
      20'h0eb73: out <= 12'h603;
      20'h0eb74: out <= 12'h603;
      20'h0eb75: out <= 12'h603;
      20'h0eb76: out <= 12'h603;
      20'h0eb77: out <= 12'h603;
      20'h0eb78: out <= 12'h603;
      20'h0eb79: out <= 12'h603;
      20'h0eb7a: out <= 12'h603;
      20'h0eb7b: out <= 12'h603;
      20'h0eb7c: out <= 12'h603;
      20'h0eb7d: out <= 12'h603;
      20'h0eb7e: out <= 12'h603;
      20'h0eb7f: out <= 12'h603;
      20'h0eb80: out <= 12'hfff;
      20'h0eb81: out <= 12'hfff;
      20'h0eb82: out <= 12'hc7f;
      20'h0eb83: out <= 12'hc7f;
      20'h0eb84: out <= 12'hc7f;
      20'h0eb85: out <= 12'hc7f;
      20'h0eb86: out <= 12'hc7f;
      20'h0eb87: out <= 12'hc7f;
      20'h0eb88: out <= 12'hc7f;
      20'h0eb89: out <= 12'hc7f;
      20'h0eb8a: out <= 12'hc7f;
      20'h0eb8b: out <= 12'hc7f;
      20'h0eb8c: out <= 12'hc7f;
      20'h0eb8d: out <= 12'hc7f;
      20'h0eb8e: out <= 12'hc7f;
      20'h0eb8f: out <= 12'hc7f;
      20'h0eb90: out <= 12'hc7f;
      20'h0eb91: out <= 12'hc7f;
      20'h0eb92: out <= 12'hc7f;
      20'h0eb93: out <= 12'hc7f;
      20'h0eb94: out <= 12'hc7f;
      20'h0eb95: out <= 12'hc7f;
      20'h0eb96: out <= 12'hc7f;
      20'h0eb97: out <= 12'hc7f;
      20'h0eb98: out <= 12'hc7f;
      20'h0eb99: out <= 12'hc7f;
      20'h0eb9a: out <= 12'hc7f;
      20'h0eb9b: out <= 12'hc7f;
      20'h0eb9c: out <= 12'hc7f;
      20'h0eb9d: out <= 12'hc7f;
      20'h0eb9e: out <= 12'hc7f;
      20'h0eb9f: out <= 12'hc7f;
      20'h0eba0: out <= 12'hc7f;
      20'h0eba1: out <= 12'hc7f;
      20'h0eba2: out <= 12'hc7f;
      20'h0eba3: out <= 12'hc7f;
      20'h0eba4: out <= 12'hc7f;
      20'h0eba5: out <= 12'hc7f;
      20'h0eba6: out <= 12'h72f;
      20'h0eba7: out <= 12'h72f;
      20'h0eba8: out <= 12'h603;
      20'h0eba9: out <= 12'h603;
      20'h0ebaa: out <= 12'h603;
      20'h0ebab: out <= 12'h603;
      20'h0ebac: out <= 12'h603;
      20'h0ebad: out <= 12'h603;
      20'h0ebae: out <= 12'h603;
      20'h0ebaf: out <= 12'h603;
      20'h0ebb0: out <= 12'h603;
      20'h0ebb1: out <= 12'h603;
      20'h0ebb2: out <= 12'h603;
      20'h0ebb3: out <= 12'h603;
      20'h0ebb4: out <= 12'h603;
      20'h0ebb5: out <= 12'h603;
      20'h0ebb6: out <= 12'h603;
      20'h0ebb7: out <= 12'h603;
      20'h0ebb8: out <= 12'h603;
      20'h0ebb9: out <= 12'h603;
      20'h0ebba: out <= 12'h603;
      20'h0ebbb: out <= 12'h603;
      20'h0ebbc: out <= 12'h603;
      20'h0ebbd: out <= 12'h603;
      20'h0ebbe: out <= 12'h603;
      20'h0ebbf: out <= 12'h603;
      20'h0ebc0: out <= 12'h603;
      20'h0ebc1: out <= 12'h603;
      20'h0ebc2: out <= 12'h603;
      20'h0ebc3: out <= 12'h603;
      20'h0ebc4: out <= 12'h603;
      20'h0ebc5: out <= 12'h603;
      20'h0ebc6: out <= 12'h603;
      20'h0ebc7: out <= 12'h603;
      20'h0ebc8: out <= 12'h603;
      20'h0ebc9: out <= 12'h603;
      20'h0ebca: out <= 12'h603;
      20'h0ebcb: out <= 12'h603;
      20'h0ebcc: out <= 12'h603;
      20'h0ebcd: out <= 12'h603;
      20'h0ebce: out <= 12'h603;
      20'h0ebcf: out <= 12'h603;
      20'h0ebd0: out <= 12'h603;
      20'h0ebd1: out <= 12'h603;
      20'h0ebd2: out <= 12'h603;
      20'h0ebd3: out <= 12'h603;
      20'h0ebd4: out <= 12'h603;
      20'h0ebd5: out <= 12'h603;
      20'h0ebd6: out <= 12'h603;
      20'h0ebd7: out <= 12'h603;
      20'h0ebd8: out <= 12'h603;
      20'h0ebd9: out <= 12'h603;
      20'h0ebda: out <= 12'h603;
      20'h0ebdb: out <= 12'h603;
      20'h0ebdc: out <= 12'h603;
      20'h0ebdd: out <= 12'h603;
      20'h0ebde: out <= 12'h603;
      20'h0ebdf: out <= 12'h603;
      20'h0ebe0: out <= 12'h603;
      20'h0ebe1: out <= 12'h603;
      20'h0ebe2: out <= 12'h603;
      20'h0ebe3: out <= 12'h603;
      20'h0ebe4: out <= 12'h603;
      20'h0ebe5: out <= 12'h603;
      20'h0ebe6: out <= 12'h603;
      20'h0ebe7: out <= 12'h603;
      20'h0ebe8: out <= 12'h603;
      20'h0ebe9: out <= 12'h603;
      20'h0ebea: out <= 12'h603;
      20'h0ebeb: out <= 12'h603;
      20'h0ebec: out <= 12'h603;
      20'h0ebed: out <= 12'h603;
      20'h0ebee: out <= 12'h603;
      20'h0ebef: out <= 12'h603;
      20'h0ebf0: out <= 12'h603;
      20'h0ebf1: out <= 12'h603;
      20'h0ebf2: out <= 12'h603;
      20'h0ebf3: out <= 12'h603;
      20'h0ebf4: out <= 12'h603;
      20'h0ebf5: out <= 12'h603;
      20'h0ebf6: out <= 12'h603;
      20'h0ebf7: out <= 12'h603;
      20'h0ebf8: out <= 12'h603;
      20'h0ebf9: out <= 12'h603;
      20'h0ebfa: out <= 12'h603;
      20'h0ebfb: out <= 12'h603;
      20'h0ebfc: out <= 12'h603;
      20'h0ebfd: out <= 12'h603;
      20'h0ebfe: out <= 12'h603;
      20'h0ebff: out <= 12'h603;
      20'h0ec00: out <= 12'hb27;
      20'h0ec01: out <= 12'hb27;
      20'h0ec02: out <= 12'hb27;
      20'h0ec03: out <= 12'hb27;
      20'h0ec04: out <= 12'hb27;
      20'h0ec05: out <= 12'hb27;
      20'h0ec06: out <= 12'hb27;
      20'h0ec07: out <= 12'hb27;
      20'h0ec08: out <= 12'h000;
      20'h0ec09: out <= 12'h000;
      20'h0ec0a: out <= 12'h000;
      20'h0ec0b: out <= 12'h000;
      20'h0ec0c: out <= 12'h000;
      20'h0ec0d: out <= 12'h000;
      20'h0ec0e: out <= 12'h000;
      20'h0ec0f: out <= 12'h000;
      20'h0ec10: out <= 12'h000;
      20'h0ec11: out <= 12'h000;
      20'h0ec12: out <= 12'h000;
      20'h0ec13: out <= 12'h000;
      20'h0ec14: out <= 12'h000;
      20'h0ec15: out <= 12'h000;
      20'h0ec16: out <= 12'h000;
      20'h0ec17: out <= 12'h000;
      20'h0ec18: out <= 12'h000;
      20'h0ec19: out <= 12'h000;
      20'h0ec1a: out <= 12'h000;
      20'h0ec1b: out <= 12'h000;
      20'h0ec1c: out <= 12'h000;
      20'h0ec1d: out <= 12'h000;
      20'h0ec1e: out <= 12'h000;
      20'h0ec1f: out <= 12'h000;
      20'h0ec20: out <= 12'h000;
      20'h0ec21: out <= 12'h000;
      20'h0ec22: out <= 12'h000;
      20'h0ec23: out <= 12'h000;
      20'h0ec24: out <= 12'h000;
      20'h0ec25: out <= 12'h000;
      20'h0ec26: out <= 12'h000;
      20'h0ec27: out <= 12'h000;
      20'h0ec28: out <= 12'h999;
      20'h0ec29: out <= 12'h999;
      20'h0ec2a: out <= 12'h999;
      20'h0ec2b: out <= 12'h999;
      20'h0ec2c: out <= 12'h999;
      20'h0ec2d: out <= 12'h999;
      20'h0ec2e: out <= 12'h999;
      20'h0ec2f: out <= 12'h999;
      20'h0ec30: out <= 12'hbbb;
      20'h0ec31: out <= 12'hbbb;
      20'h0ec32: out <= 12'hbbb;
      20'h0ec33: out <= 12'hbbb;
      20'h0ec34: out <= 12'hbbb;
      20'h0ec35: out <= 12'hbbb;
      20'h0ec36: out <= 12'hbbb;
      20'h0ec37: out <= 12'hbbb;
      20'h0ec38: out <= 12'h000;
      20'h0ec39: out <= 12'h000;
      20'h0ec3a: out <= 12'h000;
      20'h0ec3b: out <= 12'h000;
      20'h0ec3c: out <= 12'h000;
      20'h0ec3d: out <= 12'h000;
      20'h0ec3e: out <= 12'h000;
      20'h0ec3f: out <= 12'h000;
      20'h0ec40: out <= 12'hfff;
      20'h0ec41: out <= 12'hfff;
      20'h0ec42: out <= 12'hbbb;
      20'h0ec43: out <= 12'h666;
      20'h0ec44: out <= 12'h666;
      20'h0ec45: out <= 12'h666;
      20'h0ec46: out <= 12'hfff;
      20'h0ec47: out <= 12'hfff;
      20'h0ec48: out <= 12'h666;
      20'h0ec49: out <= 12'h666;
      20'h0ec4a: out <= 12'h666;
      20'h0ec4b: out <= 12'hfff;
      20'h0ec4c: out <= 12'h666;
      20'h0ec4d: out <= 12'h666;
      20'h0ec4e: out <= 12'h666;
      20'h0ec4f: out <= 12'h666;
      20'h0ec50: out <= 12'h666;
      20'h0ec51: out <= 12'h666;
      20'h0ec52: out <= 12'h666;
      20'h0ec53: out <= 12'h666;
      20'h0ec54: out <= 12'hfff;
      20'h0ec55: out <= 12'h666;
      20'h0ec56: out <= 12'h666;
      20'h0ec57: out <= 12'h666;
      20'h0ec58: out <= 12'hfff;
      20'h0ec59: out <= 12'h666;
      20'h0ec5a: out <= 12'h666;
      20'h0ec5b: out <= 12'h666;
      20'h0ec5c: out <= 12'hfff;
      20'h0ec5d: out <= 12'hfff;
      20'h0ec5e: out <= 12'hfff;
      20'h0ec5f: out <= 12'h666;
      20'h0ec60: out <= 12'h666;
      20'h0ec61: out <= 12'h666;
      20'h0ec62: out <= 12'h666;
      20'h0ec63: out <= 12'h666;
      20'h0ec64: out <= 12'hfff;
      20'h0ec65: out <= 12'hfff;
      20'h0ec66: out <= 12'h666;
      20'h0ec67: out <= 12'h666;
      20'h0ec68: out <= 12'h666;
      20'h0ec69: out <= 12'h666;
      20'h0ec6a: out <= 12'h666;
      20'h0ec6b: out <= 12'h666;
      20'h0ec6c: out <= 12'hfff;
      20'h0ec6d: out <= 12'hbbb;
      20'h0ec6e: out <= 12'h666;
      20'h0ec6f: out <= 12'h666;
      20'h0ec70: out <= 12'h603;
      20'h0ec71: out <= 12'h603;
      20'h0ec72: out <= 12'h603;
      20'h0ec73: out <= 12'h603;
      20'h0ec74: out <= 12'h603;
      20'h0ec75: out <= 12'h603;
      20'h0ec76: out <= 12'h603;
      20'h0ec77: out <= 12'h603;
      20'h0ec78: out <= 12'h603;
      20'h0ec79: out <= 12'h603;
      20'h0ec7a: out <= 12'h603;
      20'h0ec7b: out <= 12'h603;
      20'h0ec7c: out <= 12'h603;
      20'h0ec7d: out <= 12'h603;
      20'h0ec7e: out <= 12'h603;
      20'h0ec7f: out <= 12'h603;
      20'h0ec80: out <= 12'h603;
      20'h0ec81: out <= 12'h603;
      20'h0ec82: out <= 12'h603;
      20'h0ec83: out <= 12'h603;
      20'h0ec84: out <= 12'h603;
      20'h0ec85: out <= 12'h603;
      20'h0ec86: out <= 12'h603;
      20'h0ec87: out <= 12'h603;
      20'h0ec88: out <= 12'h603;
      20'h0ec89: out <= 12'h603;
      20'h0ec8a: out <= 12'h603;
      20'h0ec8b: out <= 12'h603;
      20'h0ec8c: out <= 12'h603;
      20'h0ec8d: out <= 12'h603;
      20'h0ec8e: out <= 12'h603;
      20'h0ec8f: out <= 12'h603;
      20'h0ec90: out <= 12'h603;
      20'h0ec91: out <= 12'h603;
      20'h0ec92: out <= 12'h603;
      20'h0ec93: out <= 12'h603;
      20'h0ec94: out <= 12'h603;
      20'h0ec95: out <= 12'h603;
      20'h0ec96: out <= 12'h603;
      20'h0ec97: out <= 12'h603;
      20'h0ec98: out <= 12'hfff;
      20'h0ec99: out <= 12'hfff;
      20'h0ec9a: out <= 12'hc7f;
      20'h0ec9b: out <= 12'h000;
      20'h0ec9c: out <= 12'h000;
      20'h0ec9d: out <= 12'h000;
      20'h0ec9e: out <= 12'h000;
      20'h0ec9f: out <= 12'h000;
      20'h0eca0: out <= 12'h000;
      20'h0eca1: out <= 12'h000;
      20'h0eca2: out <= 12'hc7f;
      20'h0eca3: out <= 12'hc7f;
      20'h0eca4: out <= 12'h000;
      20'h0eca5: out <= 12'h000;
      20'h0eca6: out <= 12'hc7f;
      20'h0eca7: out <= 12'hc7f;
      20'h0eca8: out <= 12'hc7f;
      20'h0eca9: out <= 12'hc7f;
      20'h0ecaa: out <= 12'h000;
      20'h0ecab: out <= 12'h000;
      20'h0ecac: out <= 12'hc7f;
      20'h0ecad: out <= 12'h000;
      20'h0ecae: out <= 12'h000;
      20'h0ecaf: out <= 12'h000;
      20'h0ecb0: out <= 12'h000;
      20'h0ecb1: out <= 12'h000;
      20'h0ecb2: out <= 12'h000;
      20'h0ecb3: out <= 12'h000;
      20'h0ecb4: out <= 12'h000;
      20'h0ecb5: out <= 12'hc7f;
      20'h0ecb6: out <= 12'h000;
      20'h0ecb7: out <= 12'h000;
      20'h0ecb8: out <= 12'h000;
      20'h0ecb9: out <= 12'h000;
      20'h0ecba: out <= 12'h000;
      20'h0ecbb: out <= 12'h000;
      20'h0ecbc: out <= 12'h000;
      20'h0ecbd: out <= 12'hc7f;
      20'h0ecbe: out <= 12'h72f;
      20'h0ecbf: out <= 12'h72f;
      20'h0ecc0: out <= 12'h603;
      20'h0ecc1: out <= 12'h603;
      20'h0ecc2: out <= 12'h603;
      20'h0ecc3: out <= 12'h603;
      20'h0ecc4: out <= 12'h603;
      20'h0ecc5: out <= 12'h603;
      20'h0ecc6: out <= 12'h603;
      20'h0ecc7: out <= 12'h603;
      20'h0ecc8: out <= 12'h603;
      20'h0ecc9: out <= 12'h603;
      20'h0ecca: out <= 12'h603;
      20'h0eccb: out <= 12'h603;
      20'h0eccc: out <= 12'h603;
      20'h0eccd: out <= 12'h603;
      20'h0ecce: out <= 12'h603;
      20'h0eccf: out <= 12'h603;
      20'h0ecd0: out <= 12'h603;
      20'h0ecd1: out <= 12'h603;
      20'h0ecd2: out <= 12'h603;
      20'h0ecd3: out <= 12'h603;
      20'h0ecd4: out <= 12'h603;
      20'h0ecd5: out <= 12'h603;
      20'h0ecd6: out <= 12'h603;
      20'h0ecd7: out <= 12'h603;
      20'h0ecd8: out <= 12'h603;
      20'h0ecd9: out <= 12'h603;
      20'h0ecda: out <= 12'h603;
      20'h0ecdb: out <= 12'h603;
      20'h0ecdc: out <= 12'h603;
      20'h0ecdd: out <= 12'h603;
      20'h0ecde: out <= 12'h603;
      20'h0ecdf: out <= 12'h603;
      20'h0ece0: out <= 12'h603;
      20'h0ece1: out <= 12'h603;
      20'h0ece2: out <= 12'h603;
      20'h0ece3: out <= 12'h603;
      20'h0ece4: out <= 12'h603;
      20'h0ece5: out <= 12'h603;
      20'h0ece6: out <= 12'h603;
      20'h0ece7: out <= 12'h603;
      20'h0ece8: out <= 12'h603;
      20'h0ece9: out <= 12'h603;
      20'h0ecea: out <= 12'h603;
      20'h0eceb: out <= 12'h603;
      20'h0ecec: out <= 12'h603;
      20'h0eced: out <= 12'h603;
      20'h0ecee: out <= 12'h603;
      20'h0ecef: out <= 12'h603;
      20'h0ecf0: out <= 12'h603;
      20'h0ecf1: out <= 12'h603;
      20'h0ecf2: out <= 12'h603;
      20'h0ecf3: out <= 12'h603;
      20'h0ecf4: out <= 12'h603;
      20'h0ecf5: out <= 12'h603;
      20'h0ecf6: out <= 12'h603;
      20'h0ecf7: out <= 12'h603;
      20'h0ecf8: out <= 12'h603;
      20'h0ecf9: out <= 12'h603;
      20'h0ecfa: out <= 12'h603;
      20'h0ecfb: out <= 12'h603;
      20'h0ecfc: out <= 12'h603;
      20'h0ecfd: out <= 12'h603;
      20'h0ecfe: out <= 12'h603;
      20'h0ecff: out <= 12'h603;
      20'h0ed00: out <= 12'h603;
      20'h0ed01: out <= 12'h603;
      20'h0ed02: out <= 12'h603;
      20'h0ed03: out <= 12'h603;
      20'h0ed04: out <= 12'h603;
      20'h0ed05: out <= 12'h603;
      20'h0ed06: out <= 12'h603;
      20'h0ed07: out <= 12'h603;
      20'h0ed08: out <= 12'h603;
      20'h0ed09: out <= 12'h603;
      20'h0ed0a: out <= 12'h603;
      20'h0ed0b: out <= 12'h603;
      20'h0ed0c: out <= 12'h603;
      20'h0ed0d: out <= 12'h603;
      20'h0ed0e: out <= 12'h603;
      20'h0ed0f: out <= 12'h603;
      20'h0ed10: out <= 12'h603;
      20'h0ed11: out <= 12'h603;
      20'h0ed12: out <= 12'h603;
      20'h0ed13: out <= 12'h603;
      20'h0ed14: out <= 12'h603;
      20'h0ed15: out <= 12'h603;
      20'h0ed16: out <= 12'h603;
      20'h0ed17: out <= 12'h603;
      20'h0ed18: out <= 12'hee9;
      20'h0ed19: out <= 12'hee9;
      20'h0ed1a: out <= 12'hee9;
      20'h0ed1b: out <= 12'hee9;
      20'h0ed1c: out <= 12'hee9;
      20'h0ed1d: out <= 12'hee9;
      20'h0ed1e: out <= 12'hee9;
      20'h0ed1f: out <= 12'hb27;
      20'h0ed20: out <= 12'hee9;
      20'h0ed21: out <= 12'hee9;
      20'h0ed22: out <= 12'hee9;
      20'h0ed23: out <= 12'hee9;
      20'h0ed24: out <= 12'hee9;
      20'h0ed25: out <= 12'hee9;
      20'h0ed26: out <= 12'hee9;
      20'h0ed27: out <= 12'hb27;
      20'h0ed28: out <= 12'hee9;
      20'h0ed29: out <= 12'hee9;
      20'h0ed2a: out <= 12'hee9;
      20'h0ed2b: out <= 12'hee9;
      20'h0ed2c: out <= 12'hee9;
      20'h0ed2d: out <= 12'hee9;
      20'h0ed2e: out <= 12'hee9;
      20'h0ed2f: out <= 12'hb27;
      20'h0ed30: out <= 12'hee9;
      20'h0ed31: out <= 12'hee9;
      20'h0ed32: out <= 12'hee9;
      20'h0ed33: out <= 12'hee9;
      20'h0ed34: out <= 12'hee9;
      20'h0ed35: out <= 12'hee9;
      20'h0ed36: out <= 12'hee9;
      20'h0ed37: out <= 12'hb27;
      20'h0ed38: out <= 12'hee9;
      20'h0ed39: out <= 12'hee9;
      20'h0ed3a: out <= 12'hee9;
      20'h0ed3b: out <= 12'hee9;
      20'h0ed3c: out <= 12'hee9;
      20'h0ed3d: out <= 12'hee9;
      20'h0ed3e: out <= 12'hee9;
      20'h0ed3f: out <= 12'hb27;
      20'h0ed40: out <= 12'hee9;
      20'h0ed41: out <= 12'hee9;
      20'h0ed42: out <= 12'hee9;
      20'h0ed43: out <= 12'hee9;
      20'h0ed44: out <= 12'hee9;
      20'h0ed45: out <= 12'hee9;
      20'h0ed46: out <= 12'hee9;
      20'h0ed47: out <= 12'hb27;
      20'h0ed48: out <= 12'hee9;
      20'h0ed49: out <= 12'hee9;
      20'h0ed4a: out <= 12'hee9;
      20'h0ed4b: out <= 12'hee9;
      20'h0ed4c: out <= 12'hee9;
      20'h0ed4d: out <= 12'hee9;
      20'h0ed4e: out <= 12'hee9;
      20'h0ed4f: out <= 12'hb27;
      20'h0ed50: out <= 12'hee9;
      20'h0ed51: out <= 12'hee9;
      20'h0ed52: out <= 12'hee9;
      20'h0ed53: out <= 12'hee9;
      20'h0ed54: out <= 12'hee9;
      20'h0ed55: out <= 12'hee9;
      20'h0ed56: out <= 12'hee9;
      20'h0ed57: out <= 12'hb27;
      20'h0ed58: out <= 12'hfff;
      20'h0ed59: out <= 12'hfff;
      20'h0ed5a: out <= 12'hbbb;
      20'h0ed5b: out <= 12'h666;
      20'h0ed5c: out <= 12'h666;
      20'h0ed5d: out <= 12'h666;
      20'h0ed5e: out <= 12'h666;
      20'h0ed5f: out <= 12'h666;
      20'h0ed60: out <= 12'h666;
      20'h0ed61: out <= 12'h666;
      20'h0ed62: out <= 12'h666;
      20'h0ed63: out <= 12'hfff;
      20'h0ed64: out <= 12'h666;
      20'h0ed65: out <= 12'h666;
      20'h0ed66: out <= 12'h666;
      20'h0ed67: out <= 12'h666;
      20'h0ed68: out <= 12'h666;
      20'h0ed69: out <= 12'h666;
      20'h0ed6a: out <= 12'h666;
      20'h0ed6b: out <= 12'h666;
      20'h0ed6c: out <= 12'hfff;
      20'h0ed6d: out <= 12'h666;
      20'h0ed6e: out <= 12'h666;
      20'h0ed6f: out <= 12'h666;
      20'h0ed70: out <= 12'hfff;
      20'h0ed71: out <= 12'h666;
      20'h0ed72: out <= 12'h666;
      20'h0ed73: out <= 12'h666;
      20'h0ed74: out <= 12'hfff;
      20'h0ed75: out <= 12'hfff;
      20'h0ed76: out <= 12'hfff;
      20'h0ed77: out <= 12'hfff;
      20'h0ed78: out <= 12'hfff;
      20'h0ed79: out <= 12'h666;
      20'h0ed7a: out <= 12'h666;
      20'h0ed7b: out <= 12'h666;
      20'h0ed7c: out <= 12'h666;
      20'h0ed7d: out <= 12'hfff;
      20'h0ed7e: out <= 12'h666;
      20'h0ed7f: out <= 12'h666;
      20'h0ed80: out <= 12'h666;
      20'h0ed81: out <= 12'hfff;
      20'h0ed82: out <= 12'hfff;
      20'h0ed83: out <= 12'hfff;
      20'h0ed84: out <= 12'hfff;
      20'h0ed85: out <= 12'hbbb;
      20'h0ed86: out <= 12'h666;
      20'h0ed87: out <= 12'h666;
      20'h0ed88: out <= 12'h603;
      20'h0ed89: out <= 12'h603;
      20'h0ed8a: out <= 12'h603;
      20'h0ed8b: out <= 12'h603;
      20'h0ed8c: out <= 12'h603;
      20'h0ed8d: out <= 12'h603;
      20'h0ed8e: out <= 12'h603;
      20'h0ed8f: out <= 12'h603;
      20'h0ed90: out <= 12'h603;
      20'h0ed91: out <= 12'h603;
      20'h0ed92: out <= 12'h603;
      20'h0ed93: out <= 12'h603;
      20'h0ed94: out <= 12'h603;
      20'h0ed95: out <= 12'h603;
      20'h0ed96: out <= 12'h603;
      20'h0ed97: out <= 12'h603;
      20'h0ed98: out <= 12'h603;
      20'h0ed99: out <= 12'h603;
      20'h0ed9a: out <= 12'h603;
      20'h0ed9b: out <= 12'h603;
      20'h0ed9c: out <= 12'h603;
      20'h0ed9d: out <= 12'h603;
      20'h0ed9e: out <= 12'h603;
      20'h0ed9f: out <= 12'h603;
      20'h0eda0: out <= 12'h603;
      20'h0eda1: out <= 12'h603;
      20'h0eda2: out <= 12'h603;
      20'h0eda3: out <= 12'h603;
      20'h0eda4: out <= 12'h603;
      20'h0eda5: out <= 12'h603;
      20'h0eda6: out <= 12'h603;
      20'h0eda7: out <= 12'h603;
      20'h0eda8: out <= 12'h603;
      20'h0eda9: out <= 12'h603;
      20'h0edaa: out <= 12'h603;
      20'h0edab: out <= 12'h603;
      20'h0edac: out <= 12'h603;
      20'h0edad: out <= 12'h603;
      20'h0edae: out <= 12'h603;
      20'h0edaf: out <= 12'h603;
      20'h0edb0: out <= 12'hfff;
      20'h0edb1: out <= 12'hfff;
      20'h0edb2: out <= 12'h000;
      20'h0edb3: out <= 12'h000;
      20'h0edb4: out <= 12'h000;
      20'h0edb5: out <= 12'hc7f;
      20'h0edb6: out <= 12'hc7f;
      20'h0edb7: out <= 12'hc7f;
      20'h0edb8: out <= 12'h000;
      20'h0edb9: out <= 12'h000;
      20'h0edba: out <= 12'h000;
      20'h0edbb: out <= 12'hc7f;
      20'h0edbc: out <= 12'h000;
      20'h0edbd: out <= 12'h000;
      20'h0edbe: out <= 12'hc7f;
      20'h0edbf: out <= 12'hc7f;
      20'h0edc0: out <= 12'hc7f;
      20'h0edc1: out <= 12'hc7f;
      20'h0edc2: out <= 12'h000;
      20'h0edc3: out <= 12'h000;
      20'h0edc4: out <= 12'hc7f;
      20'h0edc5: out <= 12'h000;
      20'h0edc6: out <= 12'h000;
      20'h0edc7: out <= 12'h000;
      20'h0edc8: out <= 12'hc7f;
      20'h0edc9: out <= 12'hc7f;
      20'h0edca: out <= 12'hc7f;
      20'h0edcb: out <= 12'hc7f;
      20'h0edcc: out <= 12'hc7f;
      20'h0edcd: out <= 12'hc7f;
      20'h0edce: out <= 12'h000;
      20'h0edcf: out <= 12'h000;
      20'h0edd0: out <= 12'h000;
      20'h0edd1: out <= 12'hc7f;
      20'h0edd2: out <= 12'hc7f;
      20'h0edd3: out <= 12'hc7f;
      20'h0edd4: out <= 12'h000;
      20'h0edd5: out <= 12'h000;
      20'h0edd6: out <= 12'h72f;
      20'h0edd7: out <= 12'h72f;
      20'h0edd8: out <= 12'h603;
      20'h0edd9: out <= 12'h603;
      20'h0edda: out <= 12'h603;
      20'h0eddb: out <= 12'h603;
      20'h0eddc: out <= 12'h603;
      20'h0eddd: out <= 12'h603;
      20'h0edde: out <= 12'h603;
      20'h0eddf: out <= 12'h603;
      20'h0ede0: out <= 12'h603;
      20'h0ede1: out <= 12'h603;
      20'h0ede2: out <= 12'h603;
      20'h0ede3: out <= 12'h603;
      20'h0ede4: out <= 12'h603;
      20'h0ede5: out <= 12'h603;
      20'h0ede6: out <= 12'h603;
      20'h0ede7: out <= 12'h603;
      20'h0ede8: out <= 12'h603;
      20'h0ede9: out <= 12'h603;
      20'h0edea: out <= 12'h603;
      20'h0edeb: out <= 12'h603;
      20'h0edec: out <= 12'h603;
      20'h0eded: out <= 12'h603;
      20'h0edee: out <= 12'h603;
      20'h0edef: out <= 12'h603;
      20'h0edf0: out <= 12'h603;
      20'h0edf1: out <= 12'h603;
      20'h0edf2: out <= 12'h603;
      20'h0edf3: out <= 12'h603;
      20'h0edf4: out <= 12'h603;
      20'h0edf5: out <= 12'h603;
      20'h0edf6: out <= 12'h603;
      20'h0edf7: out <= 12'h603;
      20'h0edf8: out <= 12'h603;
      20'h0edf9: out <= 12'h603;
      20'h0edfa: out <= 12'h603;
      20'h0edfb: out <= 12'h603;
      20'h0edfc: out <= 12'h603;
      20'h0edfd: out <= 12'h603;
      20'h0edfe: out <= 12'h603;
      20'h0edff: out <= 12'h603;
      20'h0ee00: out <= 12'h603;
      20'h0ee01: out <= 12'h603;
      20'h0ee02: out <= 12'h603;
      20'h0ee03: out <= 12'h603;
      20'h0ee04: out <= 12'h603;
      20'h0ee05: out <= 12'h603;
      20'h0ee06: out <= 12'h603;
      20'h0ee07: out <= 12'h603;
      20'h0ee08: out <= 12'h603;
      20'h0ee09: out <= 12'h603;
      20'h0ee0a: out <= 12'h603;
      20'h0ee0b: out <= 12'h603;
      20'h0ee0c: out <= 12'h603;
      20'h0ee0d: out <= 12'h603;
      20'h0ee0e: out <= 12'h603;
      20'h0ee0f: out <= 12'h603;
      20'h0ee10: out <= 12'h603;
      20'h0ee11: out <= 12'h603;
      20'h0ee12: out <= 12'h603;
      20'h0ee13: out <= 12'h603;
      20'h0ee14: out <= 12'h603;
      20'h0ee15: out <= 12'h603;
      20'h0ee16: out <= 12'h603;
      20'h0ee17: out <= 12'h603;
      20'h0ee18: out <= 12'h603;
      20'h0ee19: out <= 12'h603;
      20'h0ee1a: out <= 12'h603;
      20'h0ee1b: out <= 12'h603;
      20'h0ee1c: out <= 12'h603;
      20'h0ee1d: out <= 12'h603;
      20'h0ee1e: out <= 12'h603;
      20'h0ee1f: out <= 12'h603;
      20'h0ee20: out <= 12'h603;
      20'h0ee21: out <= 12'h603;
      20'h0ee22: out <= 12'h603;
      20'h0ee23: out <= 12'h603;
      20'h0ee24: out <= 12'h603;
      20'h0ee25: out <= 12'h603;
      20'h0ee26: out <= 12'h603;
      20'h0ee27: out <= 12'h603;
      20'h0ee28: out <= 12'h603;
      20'h0ee29: out <= 12'h603;
      20'h0ee2a: out <= 12'h603;
      20'h0ee2b: out <= 12'h603;
      20'h0ee2c: out <= 12'h603;
      20'h0ee2d: out <= 12'h603;
      20'h0ee2e: out <= 12'h603;
      20'h0ee2f: out <= 12'h603;
      20'h0ee30: out <= 12'hee9;
      20'h0ee31: out <= 12'hf87;
      20'h0ee32: out <= 12'hf87;
      20'h0ee33: out <= 12'hf87;
      20'h0ee34: out <= 12'hf87;
      20'h0ee35: out <= 12'hf87;
      20'h0ee36: out <= 12'hf87;
      20'h0ee37: out <= 12'hb27;
      20'h0ee38: out <= 12'hee9;
      20'h0ee39: out <= 12'hf87;
      20'h0ee3a: out <= 12'hf87;
      20'h0ee3b: out <= 12'hf87;
      20'h0ee3c: out <= 12'hf87;
      20'h0ee3d: out <= 12'hf87;
      20'h0ee3e: out <= 12'hf87;
      20'h0ee3f: out <= 12'hb27;
      20'h0ee40: out <= 12'hee9;
      20'h0ee41: out <= 12'hf87;
      20'h0ee42: out <= 12'hf87;
      20'h0ee43: out <= 12'hf87;
      20'h0ee44: out <= 12'hf87;
      20'h0ee45: out <= 12'hf87;
      20'h0ee46: out <= 12'hf87;
      20'h0ee47: out <= 12'hb27;
      20'h0ee48: out <= 12'hee9;
      20'h0ee49: out <= 12'hf87;
      20'h0ee4a: out <= 12'hf87;
      20'h0ee4b: out <= 12'hf87;
      20'h0ee4c: out <= 12'hf87;
      20'h0ee4d: out <= 12'hf87;
      20'h0ee4e: out <= 12'hf87;
      20'h0ee4f: out <= 12'hb27;
      20'h0ee50: out <= 12'hee9;
      20'h0ee51: out <= 12'hf87;
      20'h0ee52: out <= 12'hf87;
      20'h0ee53: out <= 12'hf87;
      20'h0ee54: out <= 12'hf87;
      20'h0ee55: out <= 12'hf87;
      20'h0ee56: out <= 12'hf87;
      20'h0ee57: out <= 12'hb27;
      20'h0ee58: out <= 12'hee9;
      20'h0ee59: out <= 12'hf87;
      20'h0ee5a: out <= 12'hf87;
      20'h0ee5b: out <= 12'hf87;
      20'h0ee5c: out <= 12'hf87;
      20'h0ee5d: out <= 12'hf87;
      20'h0ee5e: out <= 12'hf87;
      20'h0ee5f: out <= 12'hb27;
      20'h0ee60: out <= 12'hee9;
      20'h0ee61: out <= 12'hf87;
      20'h0ee62: out <= 12'hf87;
      20'h0ee63: out <= 12'hf87;
      20'h0ee64: out <= 12'hf87;
      20'h0ee65: out <= 12'hf87;
      20'h0ee66: out <= 12'hf87;
      20'h0ee67: out <= 12'hb27;
      20'h0ee68: out <= 12'hee9;
      20'h0ee69: out <= 12'hf87;
      20'h0ee6a: out <= 12'hf87;
      20'h0ee6b: out <= 12'hf87;
      20'h0ee6c: out <= 12'hf87;
      20'h0ee6d: out <= 12'hf87;
      20'h0ee6e: out <= 12'hf87;
      20'h0ee6f: out <= 12'hb27;
      20'h0ee70: out <= 12'hfff;
      20'h0ee71: out <= 12'hfff;
      20'h0ee72: out <= 12'hbbb;
      20'h0ee73: out <= 12'h666;
      20'h0ee74: out <= 12'h666;
      20'h0ee75: out <= 12'h666;
      20'h0ee76: out <= 12'h666;
      20'h0ee77: out <= 12'h666;
      20'h0ee78: out <= 12'h666;
      20'h0ee79: out <= 12'h666;
      20'h0ee7a: out <= 12'hfff;
      20'h0ee7b: out <= 12'hfff;
      20'h0ee7c: out <= 12'h666;
      20'h0ee7d: out <= 12'h666;
      20'h0ee7e: out <= 12'h666;
      20'h0ee7f: out <= 12'hfff;
      20'h0ee80: out <= 12'hfff;
      20'h0ee81: out <= 12'h666;
      20'h0ee82: out <= 12'h666;
      20'h0ee83: out <= 12'h666;
      20'h0ee84: out <= 12'hfff;
      20'h0ee85: out <= 12'h666;
      20'h0ee86: out <= 12'h666;
      20'h0ee87: out <= 12'h666;
      20'h0ee88: out <= 12'hfff;
      20'h0ee89: out <= 12'h666;
      20'h0ee8a: out <= 12'h666;
      20'h0ee8b: out <= 12'h666;
      20'h0ee8c: out <= 12'hfff;
      20'h0ee8d: out <= 12'h666;
      20'h0ee8e: out <= 12'h666;
      20'h0ee8f: out <= 12'h666;
      20'h0ee90: out <= 12'hfff;
      20'h0ee91: out <= 12'h666;
      20'h0ee92: out <= 12'h666;
      20'h0ee93: out <= 12'h666;
      20'h0ee94: out <= 12'h666;
      20'h0ee95: out <= 12'hfff;
      20'h0ee96: out <= 12'h666;
      20'h0ee97: out <= 12'h666;
      20'h0ee98: out <= 12'h666;
      20'h0ee99: out <= 12'hfff;
      20'h0ee9a: out <= 12'hfff;
      20'h0ee9b: out <= 12'hfff;
      20'h0ee9c: out <= 12'hfff;
      20'h0ee9d: out <= 12'hbbb;
      20'h0ee9e: out <= 12'h666;
      20'h0ee9f: out <= 12'h666;
      20'h0eea0: out <= 12'h603;
      20'h0eea1: out <= 12'h603;
      20'h0eea2: out <= 12'h603;
      20'h0eea3: out <= 12'h603;
      20'h0eea4: out <= 12'h603;
      20'h0eea5: out <= 12'h603;
      20'h0eea6: out <= 12'h603;
      20'h0eea7: out <= 12'h603;
      20'h0eea8: out <= 12'h603;
      20'h0eea9: out <= 12'h603;
      20'h0eeaa: out <= 12'h603;
      20'h0eeab: out <= 12'h603;
      20'h0eeac: out <= 12'h603;
      20'h0eead: out <= 12'h603;
      20'h0eeae: out <= 12'h603;
      20'h0eeaf: out <= 12'h603;
      20'h0eeb0: out <= 12'h603;
      20'h0eeb1: out <= 12'h603;
      20'h0eeb2: out <= 12'h603;
      20'h0eeb3: out <= 12'h603;
      20'h0eeb4: out <= 12'h603;
      20'h0eeb5: out <= 12'h603;
      20'h0eeb6: out <= 12'h603;
      20'h0eeb7: out <= 12'h603;
      20'h0eeb8: out <= 12'h603;
      20'h0eeb9: out <= 12'h603;
      20'h0eeba: out <= 12'h603;
      20'h0eebb: out <= 12'h603;
      20'h0eebc: out <= 12'h603;
      20'h0eebd: out <= 12'h603;
      20'h0eebe: out <= 12'h603;
      20'h0eebf: out <= 12'h603;
      20'h0eec0: out <= 12'h603;
      20'h0eec1: out <= 12'h603;
      20'h0eec2: out <= 12'h603;
      20'h0eec3: out <= 12'h603;
      20'h0eec4: out <= 12'h603;
      20'h0eec5: out <= 12'h603;
      20'h0eec6: out <= 12'h603;
      20'h0eec7: out <= 12'h603;
      20'h0eec8: out <= 12'hfff;
      20'h0eec9: out <= 12'hfff;
      20'h0eeca: out <= 12'h000;
      20'h0eecb: out <= 12'h000;
      20'h0eecc: out <= 12'h000;
      20'h0eecd: out <= 12'hc7f;
      20'h0eece: out <= 12'hc7f;
      20'h0eecf: out <= 12'hc7f;
      20'h0eed0: out <= 12'h000;
      20'h0eed1: out <= 12'h000;
      20'h0eed2: out <= 12'h000;
      20'h0eed3: out <= 12'hc7f;
      20'h0eed4: out <= 12'h000;
      20'h0eed5: out <= 12'h000;
      20'h0eed6: out <= 12'h000;
      20'h0eed7: out <= 12'hc7f;
      20'h0eed8: out <= 12'hc7f;
      20'h0eed9: out <= 12'h000;
      20'h0eeda: out <= 12'h000;
      20'h0eedb: out <= 12'h000;
      20'h0eedc: out <= 12'hc7f;
      20'h0eedd: out <= 12'h000;
      20'h0eede: out <= 12'h000;
      20'h0eedf: out <= 12'h000;
      20'h0eee0: out <= 12'h000;
      20'h0eee1: out <= 12'h000;
      20'h0eee2: out <= 12'hc7f;
      20'h0eee3: out <= 12'hc7f;
      20'h0eee4: out <= 12'hc7f;
      20'h0eee5: out <= 12'hc7f;
      20'h0eee6: out <= 12'h000;
      20'h0eee7: out <= 12'h000;
      20'h0eee8: out <= 12'h000;
      20'h0eee9: out <= 12'h000;
      20'h0eeea: out <= 12'h000;
      20'h0eeeb: out <= 12'h000;
      20'h0eeec: out <= 12'h000;
      20'h0eeed: out <= 12'hc7f;
      20'h0eeee: out <= 12'h72f;
      20'h0eeef: out <= 12'h72f;
      20'h0eef0: out <= 12'h603;
      20'h0eef1: out <= 12'h603;
      20'h0eef2: out <= 12'h603;
      20'h0eef3: out <= 12'h603;
      20'h0eef4: out <= 12'h603;
      20'h0eef5: out <= 12'h603;
      20'h0eef6: out <= 12'h603;
      20'h0eef7: out <= 12'h603;
      20'h0eef8: out <= 12'h603;
      20'h0eef9: out <= 12'h603;
      20'h0eefa: out <= 12'h603;
      20'h0eefb: out <= 12'h603;
      20'h0eefc: out <= 12'h603;
      20'h0eefd: out <= 12'h603;
      20'h0eefe: out <= 12'h603;
      20'h0eeff: out <= 12'h603;
      20'h0ef00: out <= 12'h603;
      20'h0ef01: out <= 12'h603;
      20'h0ef02: out <= 12'h603;
      20'h0ef03: out <= 12'h603;
      20'h0ef04: out <= 12'h603;
      20'h0ef05: out <= 12'h603;
      20'h0ef06: out <= 12'h603;
      20'h0ef07: out <= 12'h603;
      20'h0ef08: out <= 12'h603;
      20'h0ef09: out <= 12'h603;
      20'h0ef0a: out <= 12'h603;
      20'h0ef0b: out <= 12'h603;
      20'h0ef0c: out <= 12'h603;
      20'h0ef0d: out <= 12'h603;
      20'h0ef0e: out <= 12'h603;
      20'h0ef0f: out <= 12'h603;
      20'h0ef10: out <= 12'h603;
      20'h0ef11: out <= 12'h603;
      20'h0ef12: out <= 12'h603;
      20'h0ef13: out <= 12'h603;
      20'h0ef14: out <= 12'h603;
      20'h0ef15: out <= 12'h603;
      20'h0ef16: out <= 12'h603;
      20'h0ef17: out <= 12'h603;
      20'h0ef18: out <= 12'h603;
      20'h0ef19: out <= 12'h603;
      20'h0ef1a: out <= 12'h603;
      20'h0ef1b: out <= 12'h603;
      20'h0ef1c: out <= 12'h603;
      20'h0ef1d: out <= 12'h603;
      20'h0ef1e: out <= 12'h603;
      20'h0ef1f: out <= 12'h603;
      20'h0ef20: out <= 12'h603;
      20'h0ef21: out <= 12'h603;
      20'h0ef22: out <= 12'h603;
      20'h0ef23: out <= 12'h603;
      20'h0ef24: out <= 12'h603;
      20'h0ef25: out <= 12'h603;
      20'h0ef26: out <= 12'h603;
      20'h0ef27: out <= 12'h603;
      20'h0ef28: out <= 12'h603;
      20'h0ef29: out <= 12'h603;
      20'h0ef2a: out <= 12'h603;
      20'h0ef2b: out <= 12'h603;
      20'h0ef2c: out <= 12'h603;
      20'h0ef2d: out <= 12'h603;
      20'h0ef2e: out <= 12'h603;
      20'h0ef2f: out <= 12'h603;
      20'h0ef30: out <= 12'h603;
      20'h0ef31: out <= 12'h603;
      20'h0ef32: out <= 12'h603;
      20'h0ef33: out <= 12'h603;
      20'h0ef34: out <= 12'h603;
      20'h0ef35: out <= 12'h603;
      20'h0ef36: out <= 12'h603;
      20'h0ef37: out <= 12'h603;
      20'h0ef38: out <= 12'h603;
      20'h0ef39: out <= 12'h603;
      20'h0ef3a: out <= 12'h603;
      20'h0ef3b: out <= 12'h603;
      20'h0ef3c: out <= 12'h603;
      20'h0ef3d: out <= 12'h603;
      20'h0ef3e: out <= 12'h603;
      20'h0ef3f: out <= 12'h603;
      20'h0ef40: out <= 12'h603;
      20'h0ef41: out <= 12'h603;
      20'h0ef42: out <= 12'h603;
      20'h0ef43: out <= 12'h603;
      20'h0ef44: out <= 12'h603;
      20'h0ef45: out <= 12'h603;
      20'h0ef46: out <= 12'h603;
      20'h0ef47: out <= 12'h603;
      20'h0ef48: out <= 12'hee9;
      20'h0ef49: out <= 12'hf87;
      20'h0ef4a: out <= 12'hee9;
      20'h0ef4b: out <= 12'hee9;
      20'h0ef4c: out <= 12'hee9;
      20'h0ef4d: out <= 12'hb27;
      20'h0ef4e: out <= 12'hf87;
      20'h0ef4f: out <= 12'hb27;
      20'h0ef50: out <= 12'hee9;
      20'h0ef51: out <= 12'hf87;
      20'h0ef52: out <= 12'hee9;
      20'h0ef53: out <= 12'hee9;
      20'h0ef54: out <= 12'hee9;
      20'h0ef55: out <= 12'hb27;
      20'h0ef56: out <= 12'hf87;
      20'h0ef57: out <= 12'hb27;
      20'h0ef58: out <= 12'hee9;
      20'h0ef59: out <= 12'hf87;
      20'h0ef5a: out <= 12'hee9;
      20'h0ef5b: out <= 12'hee9;
      20'h0ef5c: out <= 12'hee9;
      20'h0ef5d: out <= 12'hb27;
      20'h0ef5e: out <= 12'hf87;
      20'h0ef5f: out <= 12'hb27;
      20'h0ef60: out <= 12'hee9;
      20'h0ef61: out <= 12'hf87;
      20'h0ef62: out <= 12'hee9;
      20'h0ef63: out <= 12'hee9;
      20'h0ef64: out <= 12'hee9;
      20'h0ef65: out <= 12'hb27;
      20'h0ef66: out <= 12'hf87;
      20'h0ef67: out <= 12'hb27;
      20'h0ef68: out <= 12'hee9;
      20'h0ef69: out <= 12'hf87;
      20'h0ef6a: out <= 12'hee9;
      20'h0ef6b: out <= 12'hee9;
      20'h0ef6c: out <= 12'hee9;
      20'h0ef6d: out <= 12'hb27;
      20'h0ef6e: out <= 12'hf87;
      20'h0ef6f: out <= 12'hb27;
      20'h0ef70: out <= 12'hee9;
      20'h0ef71: out <= 12'hf87;
      20'h0ef72: out <= 12'hee9;
      20'h0ef73: out <= 12'hee9;
      20'h0ef74: out <= 12'hee9;
      20'h0ef75: out <= 12'hb27;
      20'h0ef76: out <= 12'hf87;
      20'h0ef77: out <= 12'hb27;
      20'h0ef78: out <= 12'hee9;
      20'h0ef79: out <= 12'hf87;
      20'h0ef7a: out <= 12'hee9;
      20'h0ef7b: out <= 12'hee9;
      20'h0ef7c: out <= 12'hee9;
      20'h0ef7d: out <= 12'hb27;
      20'h0ef7e: out <= 12'hf87;
      20'h0ef7f: out <= 12'hb27;
      20'h0ef80: out <= 12'hee9;
      20'h0ef81: out <= 12'hf87;
      20'h0ef82: out <= 12'hee9;
      20'h0ef83: out <= 12'hee9;
      20'h0ef84: out <= 12'hee9;
      20'h0ef85: out <= 12'hb27;
      20'h0ef86: out <= 12'hf87;
      20'h0ef87: out <= 12'hb27;
      20'h0ef88: out <= 12'hfff;
      20'h0ef89: out <= 12'hfff;
      20'h0ef8a: out <= 12'hbbb;
      20'h0ef8b: out <= 12'h666;
      20'h0ef8c: out <= 12'h666;
      20'h0ef8d: out <= 12'h666;
      20'h0ef8e: out <= 12'hfff;
      20'h0ef8f: out <= 12'hfff;
      20'h0ef90: out <= 12'hfff;
      20'h0ef91: out <= 12'hfff;
      20'h0ef92: out <= 12'hfff;
      20'h0ef93: out <= 12'hfff;
      20'h0ef94: out <= 12'h666;
      20'h0ef95: out <= 12'h666;
      20'h0ef96: out <= 12'h666;
      20'h0ef97: out <= 12'hfff;
      20'h0ef98: out <= 12'hfff;
      20'h0ef99: out <= 12'h666;
      20'h0ef9a: out <= 12'h666;
      20'h0ef9b: out <= 12'h666;
      20'h0ef9c: out <= 12'hfff;
      20'h0ef9d: out <= 12'h666;
      20'h0ef9e: out <= 12'h666;
      20'h0ef9f: out <= 12'h666;
      20'h0efa0: out <= 12'h666;
      20'h0efa1: out <= 12'h666;
      20'h0efa2: out <= 12'h666;
      20'h0efa3: out <= 12'h666;
      20'h0efa4: out <= 12'hfff;
      20'h0efa5: out <= 12'hfff;
      20'h0efa6: out <= 12'h666;
      20'h0efa7: out <= 12'h666;
      20'h0efa8: out <= 12'h666;
      20'h0efa9: out <= 12'h666;
      20'h0efaa: out <= 12'h666;
      20'h0efab: out <= 12'h666;
      20'h0efac: out <= 12'hfff;
      20'h0efad: out <= 12'hfff;
      20'h0efae: out <= 12'h666;
      20'h0efaf: out <= 12'h666;
      20'h0efb0: out <= 12'h666;
      20'h0efb1: out <= 12'h666;
      20'h0efb2: out <= 12'h666;
      20'h0efb3: out <= 12'h666;
      20'h0efb4: out <= 12'h666;
      20'h0efb5: out <= 12'hbbb;
      20'h0efb6: out <= 12'h666;
      20'h0efb7: out <= 12'h666;
      20'h0efb8: out <= 12'h603;
      20'h0efb9: out <= 12'h603;
      20'h0efba: out <= 12'h603;
      20'h0efbb: out <= 12'h603;
      20'h0efbc: out <= 12'h603;
      20'h0efbd: out <= 12'h603;
      20'h0efbe: out <= 12'h603;
      20'h0efbf: out <= 12'h603;
      20'h0efc0: out <= 12'h603;
      20'h0efc1: out <= 12'h603;
      20'h0efc2: out <= 12'h603;
      20'h0efc3: out <= 12'h603;
      20'h0efc4: out <= 12'h603;
      20'h0efc5: out <= 12'h603;
      20'h0efc6: out <= 12'h603;
      20'h0efc7: out <= 12'h603;
      20'h0efc8: out <= 12'h603;
      20'h0efc9: out <= 12'h603;
      20'h0efca: out <= 12'h603;
      20'h0efcb: out <= 12'h603;
      20'h0efcc: out <= 12'h603;
      20'h0efcd: out <= 12'h603;
      20'h0efce: out <= 12'h603;
      20'h0efcf: out <= 12'h603;
      20'h0efd0: out <= 12'h603;
      20'h0efd1: out <= 12'h603;
      20'h0efd2: out <= 12'h603;
      20'h0efd3: out <= 12'h603;
      20'h0efd4: out <= 12'h603;
      20'h0efd5: out <= 12'h603;
      20'h0efd6: out <= 12'h603;
      20'h0efd7: out <= 12'h603;
      20'h0efd8: out <= 12'h603;
      20'h0efd9: out <= 12'h603;
      20'h0efda: out <= 12'h603;
      20'h0efdb: out <= 12'h603;
      20'h0efdc: out <= 12'h603;
      20'h0efdd: out <= 12'h603;
      20'h0efde: out <= 12'h603;
      20'h0efdf: out <= 12'h603;
      20'h0efe0: out <= 12'hfff;
      20'h0efe1: out <= 12'hfff;
      20'h0efe2: out <= 12'h000;
      20'h0efe3: out <= 12'h000;
      20'h0efe4: out <= 12'h000;
      20'h0efe5: out <= 12'hc7f;
      20'h0efe6: out <= 12'hc7f;
      20'h0efe7: out <= 12'hc7f;
      20'h0efe8: out <= 12'h000;
      20'h0efe9: out <= 12'h000;
      20'h0efea: out <= 12'h000;
      20'h0efeb: out <= 12'hc7f;
      20'h0efec: out <= 12'hc7f;
      20'h0efed: out <= 12'h000;
      20'h0efee: out <= 12'h000;
      20'h0efef: out <= 12'hc7f;
      20'h0eff0: out <= 12'hc7f;
      20'h0eff1: out <= 12'h000;
      20'h0eff2: out <= 12'h000;
      20'h0eff3: out <= 12'hc7f;
      20'h0eff4: out <= 12'hc7f;
      20'h0eff5: out <= 12'h000;
      20'h0eff6: out <= 12'h000;
      20'h0eff7: out <= 12'h000;
      20'h0eff8: out <= 12'hc7f;
      20'h0eff9: out <= 12'hc7f;
      20'h0effa: out <= 12'hc7f;
      20'h0effb: out <= 12'hc7f;
      20'h0effc: out <= 12'hc7f;
      20'h0effd: out <= 12'hc7f;
      20'h0effe: out <= 12'h000;
      20'h0efff: out <= 12'h000;
      20'h0f000: out <= 12'h000;
      20'h0f001: out <= 12'hc7f;
      20'h0f002: out <= 12'h000;
      20'h0f003: out <= 12'h000;
      20'h0f004: out <= 12'hc7f;
      20'h0f005: out <= 12'hc7f;
      20'h0f006: out <= 12'h72f;
      20'h0f007: out <= 12'h72f;
      20'h0f008: out <= 12'h603;
      20'h0f009: out <= 12'h603;
      20'h0f00a: out <= 12'h603;
      20'h0f00b: out <= 12'h603;
      20'h0f00c: out <= 12'h603;
      20'h0f00d: out <= 12'h603;
      20'h0f00e: out <= 12'h603;
      20'h0f00f: out <= 12'h603;
      20'h0f010: out <= 12'h603;
      20'h0f011: out <= 12'h603;
      20'h0f012: out <= 12'h603;
      20'h0f013: out <= 12'h603;
      20'h0f014: out <= 12'h603;
      20'h0f015: out <= 12'h603;
      20'h0f016: out <= 12'h603;
      20'h0f017: out <= 12'h603;
      20'h0f018: out <= 12'h603;
      20'h0f019: out <= 12'h603;
      20'h0f01a: out <= 12'h603;
      20'h0f01b: out <= 12'h603;
      20'h0f01c: out <= 12'h603;
      20'h0f01d: out <= 12'h603;
      20'h0f01e: out <= 12'h603;
      20'h0f01f: out <= 12'h603;
      20'h0f020: out <= 12'h603;
      20'h0f021: out <= 12'h603;
      20'h0f022: out <= 12'h603;
      20'h0f023: out <= 12'h603;
      20'h0f024: out <= 12'h603;
      20'h0f025: out <= 12'h603;
      20'h0f026: out <= 12'h603;
      20'h0f027: out <= 12'h603;
      20'h0f028: out <= 12'h603;
      20'h0f029: out <= 12'h603;
      20'h0f02a: out <= 12'h603;
      20'h0f02b: out <= 12'h603;
      20'h0f02c: out <= 12'h603;
      20'h0f02d: out <= 12'h603;
      20'h0f02e: out <= 12'h603;
      20'h0f02f: out <= 12'h603;
      20'h0f030: out <= 12'h603;
      20'h0f031: out <= 12'h603;
      20'h0f032: out <= 12'h603;
      20'h0f033: out <= 12'h603;
      20'h0f034: out <= 12'h603;
      20'h0f035: out <= 12'h603;
      20'h0f036: out <= 12'h603;
      20'h0f037: out <= 12'h603;
      20'h0f038: out <= 12'h603;
      20'h0f039: out <= 12'h603;
      20'h0f03a: out <= 12'h603;
      20'h0f03b: out <= 12'h603;
      20'h0f03c: out <= 12'h603;
      20'h0f03d: out <= 12'h603;
      20'h0f03e: out <= 12'h603;
      20'h0f03f: out <= 12'h603;
      20'h0f040: out <= 12'h603;
      20'h0f041: out <= 12'h603;
      20'h0f042: out <= 12'h603;
      20'h0f043: out <= 12'h603;
      20'h0f044: out <= 12'h603;
      20'h0f045: out <= 12'h603;
      20'h0f046: out <= 12'h603;
      20'h0f047: out <= 12'h603;
      20'h0f048: out <= 12'h603;
      20'h0f049: out <= 12'h603;
      20'h0f04a: out <= 12'h603;
      20'h0f04b: out <= 12'h603;
      20'h0f04c: out <= 12'h603;
      20'h0f04d: out <= 12'h603;
      20'h0f04e: out <= 12'h603;
      20'h0f04f: out <= 12'h603;
      20'h0f050: out <= 12'h603;
      20'h0f051: out <= 12'h603;
      20'h0f052: out <= 12'h603;
      20'h0f053: out <= 12'h603;
      20'h0f054: out <= 12'h603;
      20'h0f055: out <= 12'h603;
      20'h0f056: out <= 12'h603;
      20'h0f057: out <= 12'h603;
      20'h0f058: out <= 12'h603;
      20'h0f059: out <= 12'h603;
      20'h0f05a: out <= 12'h603;
      20'h0f05b: out <= 12'h603;
      20'h0f05c: out <= 12'h603;
      20'h0f05d: out <= 12'h603;
      20'h0f05e: out <= 12'h603;
      20'h0f05f: out <= 12'h603;
      20'h0f060: out <= 12'hee9;
      20'h0f061: out <= 12'hf87;
      20'h0f062: out <= 12'hee9;
      20'h0f063: out <= 12'hf87;
      20'h0f064: out <= 12'hf87;
      20'h0f065: out <= 12'hb27;
      20'h0f066: out <= 12'hf87;
      20'h0f067: out <= 12'hb27;
      20'h0f068: out <= 12'hee9;
      20'h0f069: out <= 12'hf87;
      20'h0f06a: out <= 12'hee9;
      20'h0f06b: out <= 12'hf87;
      20'h0f06c: out <= 12'hf87;
      20'h0f06d: out <= 12'hb27;
      20'h0f06e: out <= 12'hf87;
      20'h0f06f: out <= 12'hb27;
      20'h0f070: out <= 12'hee9;
      20'h0f071: out <= 12'hf87;
      20'h0f072: out <= 12'hee9;
      20'h0f073: out <= 12'hf87;
      20'h0f074: out <= 12'hf87;
      20'h0f075: out <= 12'hb27;
      20'h0f076: out <= 12'hf87;
      20'h0f077: out <= 12'hb27;
      20'h0f078: out <= 12'hee9;
      20'h0f079: out <= 12'hf87;
      20'h0f07a: out <= 12'hee9;
      20'h0f07b: out <= 12'hf87;
      20'h0f07c: out <= 12'hf87;
      20'h0f07d: out <= 12'hb27;
      20'h0f07e: out <= 12'hf87;
      20'h0f07f: out <= 12'hb27;
      20'h0f080: out <= 12'hee9;
      20'h0f081: out <= 12'hf87;
      20'h0f082: out <= 12'hee9;
      20'h0f083: out <= 12'hf87;
      20'h0f084: out <= 12'hf87;
      20'h0f085: out <= 12'hb27;
      20'h0f086: out <= 12'hf87;
      20'h0f087: out <= 12'hb27;
      20'h0f088: out <= 12'hee9;
      20'h0f089: out <= 12'hf87;
      20'h0f08a: out <= 12'hee9;
      20'h0f08b: out <= 12'hf87;
      20'h0f08c: out <= 12'hf87;
      20'h0f08d: out <= 12'hb27;
      20'h0f08e: out <= 12'hf87;
      20'h0f08f: out <= 12'hb27;
      20'h0f090: out <= 12'hee9;
      20'h0f091: out <= 12'hf87;
      20'h0f092: out <= 12'hee9;
      20'h0f093: out <= 12'hf87;
      20'h0f094: out <= 12'hf87;
      20'h0f095: out <= 12'hb27;
      20'h0f096: out <= 12'hf87;
      20'h0f097: out <= 12'hb27;
      20'h0f098: out <= 12'hee9;
      20'h0f099: out <= 12'hf87;
      20'h0f09a: out <= 12'hee9;
      20'h0f09b: out <= 12'hf87;
      20'h0f09c: out <= 12'hf87;
      20'h0f09d: out <= 12'hb27;
      20'h0f09e: out <= 12'hf87;
      20'h0f09f: out <= 12'hb27;
      20'h0f0a0: out <= 12'hfff;
      20'h0f0a1: out <= 12'hfff;
      20'h0f0a2: out <= 12'hbbb;
      20'h0f0a3: out <= 12'h666;
      20'h0f0a4: out <= 12'h666;
      20'h0f0a5: out <= 12'h666;
      20'h0f0a6: out <= 12'hfff;
      20'h0f0a7: out <= 12'hfff;
      20'h0f0a8: out <= 12'hfff;
      20'h0f0a9: out <= 12'hfff;
      20'h0f0aa: out <= 12'hfff;
      20'h0f0ab: out <= 12'hfff;
      20'h0f0ac: out <= 12'h666;
      20'h0f0ad: out <= 12'h666;
      20'h0f0ae: out <= 12'h666;
      20'h0f0af: out <= 12'hfff;
      20'h0f0b0: out <= 12'hfff;
      20'h0f0b1: out <= 12'h666;
      20'h0f0b2: out <= 12'h666;
      20'h0f0b3: out <= 12'h666;
      20'h0f0b4: out <= 12'hfff;
      20'h0f0b5: out <= 12'hfff;
      20'h0f0b6: out <= 12'h666;
      20'h0f0b7: out <= 12'h666;
      20'h0f0b8: out <= 12'h666;
      20'h0f0b9: out <= 12'h666;
      20'h0f0ba: out <= 12'h666;
      20'h0f0bb: out <= 12'hfff;
      20'h0f0bc: out <= 12'hfff;
      20'h0f0bd: out <= 12'hfff;
      20'h0f0be: out <= 12'hfff;
      20'h0f0bf: out <= 12'h666;
      20'h0f0c0: out <= 12'h666;
      20'h0f0c1: out <= 12'h666;
      20'h0f0c2: out <= 12'h666;
      20'h0f0c3: out <= 12'hfff;
      20'h0f0c4: out <= 12'hfff;
      20'h0f0c5: out <= 12'hfff;
      20'h0f0c6: out <= 12'h666;
      20'h0f0c7: out <= 12'h666;
      20'h0f0c8: out <= 12'h666;
      20'h0f0c9: out <= 12'h666;
      20'h0f0ca: out <= 12'h666;
      20'h0f0cb: out <= 12'h666;
      20'h0f0cc: out <= 12'h666;
      20'h0f0cd: out <= 12'hbbb;
      20'h0f0ce: out <= 12'h666;
      20'h0f0cf: out <= 12'h666;
      20'h0f0d0: out <= 12'h603;
      20'h0f0d1: out <= 12'h603;
      20'h0f0d2: out <= 12'h603;
      20'h0f0d3: out <= 12'h603;
      20'h0f0d4: out <= 12'h603;
      20'h0f0d5: out <= 12'h603;
      20'h0f0d6: out <= 12'h603;
      20'h0f0d7: out <= 12'h603;
      20'h0f0d8: out <= 12'h603;
      20'h0f0d9: out <= 12'h603;
      20'h0f0da: out <= 12'h603;
      20'h0f0db: out <= 12'h603;
      20'h0f0dc: out <= 12'h603;
      20'h0f0dd: out <= 12'h603;
      20'h0f0de: out <= 12'h603;
      20'h0f0df: out <= 12'h603;
      20'h0f0e0: out <= 12'h603;
      20'h0f0e1: out <= 12'h603;
      20'h0f0e2: out <= 12'h603;
      20'h0f0e3: out <= 12'h603;
      20'h0f0e4: out <= 12'h603;
      20'h0f0e5: out <= 12'h603;
      20'h0f0e6: out <= 12'h603;
      20'h0f0e7: out <= 12'h603;
      20'h0f0e8: out <= 12'h603;
      20'h0f0e9: out <= 12'h603;
      20'h0f0ea: out <= 12'h603;
      20'h0f0eb: out <= 12'h603;
      20'h0f0ec: out <= 12'h603;
      20'h0f0ed: out <= 12'h603;
      20'h0f0ee: out <= 12'h603;
      20'h0f0ef: out <= 12'h603;
      20'h0f0f0: out <= 12'h603;
      20'h0f0f1: out <= 12'h603;
      20'h0f0f2: out <= 12'h603;
      20'h0f0f3: out <= 12'h603;
      20'h0f0f4: out <= 12'h603;
      20'h0f0f5: out <= 12'h603;
      20'h0f0f6: out <= 12'h603;
      20'h0f0f7: out <= 12'h603;
      20'h0f0f8: out <= 12'hfff;
      20'h0f0f9: out <= 12'hfff;
      20'h0f0fa: out <= 12'h000;
      20'h0f0fb: out <= 12'h000;
      20'h0f0fc: out <= 12'h000;
      20'h0f0fd: out <= 12'hc7f;
      20'h0f0fe: out <= 12'hc7f;
      20'h0f0ff: out <= 12'hc7f;
      20'h0f100: out <= 12'h000;
      20'h0f101: out <= 12'h000;
      20'h0f102: out <= 12'h000;
      20'h0f103: out <= 12'hc7f;
      20'h0f104: out <= 12'hc7f;
      20'h0f105: out <= 12'h000;
      20'h0f106: out <= 12'h000;
      20'h0f107: out <= 12'h000;
      20'h0f108: out <= 12'h000;
      20'h0f109: out <= 12'h000;
      20'h0f10a: out <= 12'h000;
      20'h0f10b: out <= 12'hc7f;
      20'h0f10c: out <= 12'hc7f;
      20'h0f10d: out <= 12'h000;
      20'h0f10e: out <= 12'h000;
      20'h0f10f: out <= 12'h000;
      20'h0f110: out <= 12'hc7f;
      20'h0f111: out <= 12'hc7f;
      20'h0f112: out <= 12'hc7f;
      20'h0f113: out <= 12'hc7f;
      20'h0f114: out <= 12'hc7f;
      20'h0f115: out <= 12'hc7f;
      20'h0f116: out <= 12'h000;
      20'h0f117: out <= 12'h000;
      20'h0f118: out <= 12'h000;
      20'h0f119: out <= 12'hc7f;
      20'h0f11a: out <= 12'hc7f;
      20'h0f11b: out <= 12'h000;
      20'h0f11c: out <= 12'h000;
      20'h0f11d: out <= 12'hc7f;
      20'h0f11e: out <= 12'h72f;
      20'h0f11f: out <= 12'h72f;
      20'h0f120: out <= 12'h603;
      20'h0f121: out <= 12'h603;
      20'h0f122: out <= 12'h603;
      20'h0f123: out <= 12'h603;
      20'h0f124: out <= 12'h603;
      20'h0f125: out <= 12'h603;
      20'h0f126: out <= 12'h603;
      20'h0f127: out <= 12'h603;
      20'h0f128: out <= 12'h603;
      20'h0f129: out <= 12'h603;
      20'h0f12a: out <= 12'h603;
      20'h0f12b: out <= 12'h603;
      20'h0f12c: out <= 12'h603;
      20'h0f12d: out <= 12'h603;
      20'h0f12e: out <= 12'h603;
      20'h0f12f: out <= 12'h603;
      20'h0f130: out <= 12'h603;
      20'h0f131: out <= 12'h603;
      20'h0f132: out <= 12'h603;
      20'h0f133: out <= 12'h603;
      20'h0f134: out <= 12'h603;
      20'h0f135: out <= 12'h603;
      20'h0f136: out <= 12'h603;
      20'h0f137: out <= 12'h603;
      20'h0f138: out <= 12'h603;
      20'h0f139: out <= 12'h603;
      20'h0f13a: out <= 12'h603;
      20'h0f13b: out <= 12'h603;
      20'h0f13c: out <= 12'h603;
      20'h0f13d: out <= 12'h603;
      20'h0f13e: out <= 12'h603;
      20'h0f13f: out <= 12'h603;
      20'h0f140: out <= 12'h603;
      20'h0f141: out <= 12'h603;
      20'h0f142: out <= 12'h603;
      20'h0f143: out <= 12'h603;
      20'h0f144: out <= 12'h603;
      20'h0f145: out <= 12'h603;
      20'h0f146: out <= 12'h603;
      20'h0f147: out <= 12'h603;
      20'h0f148: out <= 12'h603;
      20'h0f149: out <= 12'h603;
      20'h0f14a: out <= 12'h603;
      20'h0f14b: out <= 12'h603;
      20'h0f14c: out <= 12'h603;
      20'h0f14d: out <= 12'h603;
      20'h0f14e: out <= 12'h603;
      20'h0f14f: out <= 12'h603;
      20'h0f150: out <= 12'h603;
      20'h0f151: out <= 12'h603;
      20'h0f152: out <= 12'h603;
      20'h0f153: out <= 12'h603;
      20'h0f154: out <= 12'h603;
      20'h0f155: out <= 12'h603;
      20'h0f156: out <= 12'h603;
      20'h0f157: out <= 12'h603;
      20'h0f158: out <= 12'h603;
      20'h0f159: out <= 12'h603;
      20'h0f15a: out <= 12'h603;
      20'h0f15b: out <= 12'h603;
      20'h0f15c: out <= 12'h603;
      20'h0f15d: out <= 12'h603;
      20'h0f15e: out <= 12'h603;
      20'h0f15f: out <= 12'h603;
      20'h0f160: out <= 12'h603;
      20'h0f161: out <= 12'h603;
      20'h0f162: out <= 12'h603;
      20'h0f163: out <= 12'h603;
      20'h0f164: out <= 12'h603;
      20'h0f165: out <= 12'h603;
      20'h0f166: out <= 12'h603;
      20'h0f167: out <= 12'h603;
      20'h0f168: out <= 12'h603;
      20'h0f169: out <= 12'h603;
      20'h0f16a: out <= 12'h603;
      20'h0f16b: out <= 12'h603;
      20'h0f16c: out <= 12'h603;
      20'h0f16d: out <= 12'h603;
      20'h0f16e: out <= 12'h603;
      20'h0f16f: out <= 12'h603;
      20'h0f170: out <= 12'h603;
      20'h0f171: out <= 12'h603;
      20'h0f172: out <= 12'h603;
      20'h0f173: out <= 12'h603;
      20'h0f174: out <= 12'h603;
      20'h0f175: out <= 12'h603;
      20'h0f176: out <= 12'h603;
      20'h0f177: out <= 12'h603;
      20'h0f178: out <= 12'hee9;
      20'h0f179: out <= 12'hf87;
      20'h0f17a: out <= 12'hee9;
      20'h0f17b: out <= 12'hf87;
      20'h0f17c: out <= 12'hf87;
      20'h0f17d: out <= 12'hb27;
      20'h0f17e: out <= 12'hf87;
      20'h0f17f: out <= 12'hb27;
      20'h0f180: out <= 12'hee9;
      20'h0f181: out <= 12'hf87;
      20'h0f182: out <= 12'hee9;
      20'h0f183: out <= 12'hf87;
      20'h0f184: out <= 12'hf87;
      20'h0f185: out <= 12'hb27;
      20'h0f186: out <= 12'hf87;
      20'h0f187: out <= 12'hb27;
      20'h0f188: out <= 12'hee9;
      20'h0f189: out <= 12'hf87;
      20'h0f18a: out <= 12'hee9;
      20'h0f18b: out <= 12'hf87;
      20'h0f18c: out <= 12'hf87;
      20'h0f18d: out <= 12'hb27;
      20'h0f18e: out <= 12'hf87;
      20'h0f18f: out <= 12'hb27;
      20'h0f190: out <= 12'hee9;
      20'h0f191: out <= 12'hf87;
      20'h0f192: out <= 12'hee9;
      20'h0f193: out <= 12'hf87;
      20'h0f194: out <= 12'hf87;
      20'h0f195: out <= 12'hb27;
      20'h0f196: out <= 12'hf87;
      20'h0f197: out <= 12'hb27;
      20'h0f198: out <= 12'hee9;
      20'h0f199: out <= 12'hf87;
      20'h0f19a: out <= 12'hee9;
      20'h0f19b: out <= 12'hf87;
      20'h0f19c: out <= 12'hf87;
      20'h0f19d: out <= 12'hb27;
      20'h0f19e: out <= 12'hf87;
      20'h0f19f: out <= 12'hb27;
      20'h0f1a0: out <= 12'hee9;
      20'h0f1a1: out <= 12'hf87;
      20'h0f1a2: out <= 12'hee9;
      20'h0f1a3: out <= 12'hf87;
      20'h0f1a4: out <= 12'hf87;
      20'h0f1a5: out <= 12'hb27;
      20'h0f1a6: out <= 12'hf87;
      20'h0f1a7: out <= 12'hb27;
      20'h0f1a8: out <= 12'hee9;
      20'h0f1a9: out <= 12'hf87;
      20'h0f1aa: out <= 12'hee9;
      20'h0f1ab: out <= 12'hf87;
      20'h0f1ac: out <= 12'hf87;
      20'h0f1ad: out <= 12'hb27;
      20'h0f1ae: out <= 12'hf87;
      20'h0f1af: out <= 12'hb27;
      20'h0f1b0: out <= 12'hee9;
      20'h0f1b1: out <= 12'hf87;
      20'h0f1b2: out <= 12'hee9;
      20'h0f1b3: out <= 12'hf87;
      20'h0f1b4: out <= 12'hf87;
      20'h0f1b5: out <= 12'hb27;
      20'h0f1b6: out <= 12'hf87;
      20'h0f1b7: out <= 12'hb27;
      20'h0f1b8: out <= 12'hfff;
      20'h0f1b9: out <= 12'hfff;
      20'h0f1ba: out <= 12'hbbb;
      20'h0f1bb: out <= 12'hbbb;
      20'h0f1bc: out <= 12'hbbb;
      20'h0f1bd: out <= 12'hbbb;
      20'h0f1be: out <= 12'hbbb;
      20'h0f1bf: out <= 12'hbbb;
      20'h0f1c0: out <= 12'hbbb;
      20'h0f1c1: out <= 12'hbbb;
      20'h0f1c2: out <= 12'hbbb;
      20'h0f1c3: out <= 12'hbbb;
      20'h0f1c4: out <= 12'hbbb;
      20'h0f1c5: out <= 12'hbbb;
      20'h0f1c6: out <= 12'hbbb;
      20'h0f1c7: out <= 12'hbbb;
      20'h0f1c8: out <= 12'hbbb;
      20'h0f1c9: out <= 12'hbbb;
      20'h0f1ca: out <= 12'hbbb;
      20'h0f1cb: out <= 12'hbbb;
      20'h0f1cc: out <= 12'hbbb;
      20'h0f1cd: out <= 12'hbbb;
      20'h0f1ce: out <= 12'hbbb;
      20'h0f1cf: out <= 12'hbbb;
      20'h0f1d0: out <= 12'hbbb;
      20'h0f1d1: out <= 12'hbbb;
      20'h0f1d2: out <= 12'hbbb;
      20'h0f1d3: out <= 12'hbbb;
      20'h0f1d4: out <= 12'hbbb;
      20'h0f1d5: out <= 12'hbbb;
      20'h0f1d6: out <= 12'hbbb;
      20'h0f1d7: out <= 12'hbbb;
      20'h0f1d8: out <= 12'hbbb;
      20'h0f1d9: out <= 12'hbbb;
      20'h0f1da: out <= 12'hbbb;
      20'h0f1db: out <= 12'hbbb;
      20'h0f1dc: out <= 12'hbbb;
      20'h0f1dd: out <= 12'hbbb;
      20'h0f1de: out <= 12'hbbb;
      20'h0f1df: out <= 12'hbbb;
      20'h0f1e0: out <= 12'hbbb;
      20'h0f1e1: out <= 12'hbbb;
      20'h0f1e2: out <= 12'hbbb;
      20'h0f1e3: out <= 12'hbbb;
      20'h0f1e4: out <= 12'hbbb;
      20'h0f1e5: out <= 12'hbbb;
      20'h0f1e6: out <= 12'h666;
      20'h0f1e7: out <= 12'h666;
      20'h0f1e8: out <= 12'h603;
      20'h0f1e9: out <= 12'h603;
      20'h0f1ea: out <= 12'h603;
      20'h0f1eb: out <= 12'h603;
      20'h0f1ec: out <= 12'h603;
      20'h0f1ed: out <= 12'h603;
      20'h0f1ee: out <= 12'h603;
      20'h0f1ef: out <= 12'h603;
      20'h0f1f0: out <= 12'h603;
      20'h0f1f1: out <= 12'h603;
      20'h0f1f2: out <= 12'h603;
      20'h0f1f3: out <= 12'h603;
      20'h0f1f4: out <= 12'h603;
      20'h0f1f5: out <= 12'h603;
      20'h0f1f6: out <= 12'h603;
      20'h0f1f7: out <= 12'h603;
      20'h0f1f8: out <= 12'h603;
      20'h0f1f9: out <= 12'h603;
      20'h0f1fa: out <= 12'h603;
      20'h0f1fb: out <= 12'h603;
      20'h0f1fc: out <= 12'h603;
      20'h0f1fd: out <= 12'h603;
      20'h0f1fe: out <= 12'h603;
      20'h0f1ff: out <= 12'h603;
      20'h0f200: out <= 12'h603;
      20'h0f201: out <= 12'h603;
      20'h0f202: out <= 12'h603;
      20'h0f203: out <= 12'h603;
      20'h0f204: out <= 12'h603;
      20'h0f205: out <= 12'h603;
      20'h0f206: out <= 12'h603;
      20'h0f207: out <= 12'h603;
      20'h0f208: out <= 12'h603;
      20'h0f209: out <= 12'h603;
      20'h0f20a: out <= 12'h603;
      20'h0f20b: out <= 12'h603;
      20'h0f20c: out <= 12'h603;
      20'h0f20d: out <= 12'h603;
      20'h0f20e: out <= 12'h603;
      20'h0f20f: out <= 12'h603;
      20'h0f210: out <= 12'hfff;
      20'h0f211: out <= 12'hfff;
      20'h0f212: out <= 12'hc7f;
      20'h0f213: out <= 12'h000;
      20'h0f214: out <= 12'h000;
      20'h0f215: out <= 12'h000;
      20'h0f216: out <= 12'h000;
      20'h0f217: out <= 12'h000;
      20'h0f218: out <= 12'h000;
      20'h0f219: out <= 12'h000;
      20'h0f21a: out <= 12'hc7f;
      20'h0f21b: out <= 12'hc7f;
      20'h0f21c: out <= 12'hc7f;
      20'h0f21d: out <= 12'hc7f;
      20'h0f21e: out <= 12'h000;
      20'h0f21f: out <= 12'h000;
      20'h0f220: out <= 12'h000;
      20'h0f221: out <= 12'h000;
      20'h0f222: out <= 12'hc7f;
      20'h0f223: out <= 12'hc7f;
      20'h0f224: out <= 12'hc7f;
      20'h0f225: out <= 12'h000;
      20'h0f226: out <= 12'h000;
      20'h0f227: out <= 12'h000;
      20'h0f228: out <= 12'h000;
      20'h0f229: out <= 12'h000;
      20'h0f22a: out <= 12'h000;
      20'h0f22b: out <= 12'h000;
      20'h0f22c: out <= 12'h000;
      20'h0f22d: out <= 12'hc7f;
      20'h0f22e: out <= 12'h000;
      20'h0f22f: out <= 12'h000;
      20'h0f230: out <= 12'h000;
      20'h0f231: out <= 12'hc7f;
      20'h0f232: out <= 12'hc7f;
      20'h0f233: out <= 12'hc7f;
      20'h0f234: out <= 12'h000;
      20'h0f235: out <= 12'h000;
      20'h0f236: out <= 12'h72f;
      20'h0f237: out <= 12'h72f;
      20'h0f238: out <= 12'h603;
      20'h0f239: out <= 12'h603;
      20'h0f23a: out <= 12'h603;
      20'h0f23b: out <= 12'h603;
      20'h0f23c: out <= 12'h603;
      20'h0f23d: out <= 12'h603;
      20'h0f23e: out <= 12'h603;
      20'h0f23f: out <= 12'h603;
      20'h0f240: out <= 12'h603;
      20'h0f241: out <= 12'h603;
      20'h0f242: out <= 12'h603;
      20'h0f243: out <= 12'h603;
      20'h0f244: out <= 12'h603;
      20'h0f245: out <= 12'h603;
      20'h0f246: out <= 12'h603;
      20'h0f247: out <= 12'h603;
      20'h0f248: out <= 12'h603;
      20'h0f249: out <= 12'h603;
      20'h0f24a: out <= 12'h603;
      20'h0f24b: out <= 12'h603;
      20'h0f24c: out <= 12'h603;
      20'h0f24d: out <= 12'h603;
      20'h0f24e: out <= 12'h603;
      20'h0f24f: out <= 12'h603;
      20'h0f250: out <= 12'h603;
      20'h0f251: out <= 12'h603;
      20'h0f252: out <= 12'h603;
      20'h0f253: out <= 12'h603;
      20'h0f254: out <= 12'h603;
      20'h0f255: out <= 12'h603;
      20'h0f256: out <= 12'h603;
      20'h0f257: out <= 12'h603;
      20'h0f258: out <= 12'h603;
      20'h0f259: out <= 12'h603;
      20'h0f25a: out <= 12'h603;
      20'h0f25b: out <= 12'h603;
      20'h0f25c: out <= 12'h603;
      20'h0f25d: out <= 12'h603;
      20'h0f25e: out <= 12'h603;
      20'h0f25f: out <= 12'h603;
      20'h0f260: out <= 12'h603;
      20'h0f261: out <= 12'h603;
      20'h0f262: out <= 12'h603;
      20'h0f263: out <= 12'h603;
      20'h0f264: out <= 12'h603;
      20'h0f265: out <= 12'h603;
      20'h0f266: out <= 12'h603;
      20'h0f267: out <= 12'h603;
      20'h0f268: out <= 12'h603;
      20'h0f269: out <= 12'h603;
      20'h0f26a: out <= 12'h603;
      20'h0f26b: out <= 12'h603;
      20'h0f26c: out <= 12'h603;
      20'h0f26d: out <= 12'h603;
      20'h0f26e: out <= 12'h603;
      20'h0f26f: out <= 12'h603;
      20'h0f270: out <= 12'h603;
      20'h0f271: out <= 12'h603;
      20'h0f272: out <= 12'h603;
      20'h0f273: out <= 12'h603;
      20'h0f274: out <= 12'h603;
      20'h0f275: out <= 12'h603;
      20'h0f276: out <= 12'h603;
      20'h0f277: out <= 12'h603;
      20'h0f278: out <= 12'h603;
      20'h0f279: out <= 12'h603;
      20'h0f27a: out <= 12'h603;
      20'h0f27b: out <= 12'h603;
      20'h0f27c: out <= 12'h603;
      20'h0f27d: out <= 12'h603;
      20'h0f27e: out <= 12'h603;
      20'h0f27f: out <= 12'h603;
      20'h0f280: out <= 12'h603;
      20'h0f281: out <= 12'h603;
      20'h0f282: out <= 12'h603;
      20'h0f283: out <= 12'h603;
      20'h0f284: out <= 12'h603;
      20'h0f285: out <= 12'h603;
      20'h0f286: out <= 12'h603;
      20'h0f287: out <= 12'h603;
      20'h0f288: out <= 12'h603;
      20'h0f289: out <= 12'h603;
      20'h0f28a: out <= 12'h603;
      20'h0f28b: out <= 12'h603;
      20'h0f28c: out <= 12'h603;
      20'h0f28d: out <= 12'h603;
      20'h0f28e: out <= 12'h603;
      20'h0f28f: out <= 12'h603;
      20'h0f290: out <= 12'hee9;
      20'h0f291: out <= 12'hf87;
      20'h0f292: out <= 12'hee9;
      20'h0f293: out <= 12'hb27;
      20'h0f294: out <= 12'hb27;
      20'h0f295: out <= 12'hb27;
      20'h0f296: out <= 12'hf87;
      20'h0f297: out <= 12'hb27;
      20'h0f298: out <= 12'hee9;
      20'h0f299: out <= 12'hf87;
      20'h0f29a: out <= 12'hee9;
      20'h0f29b: out <= 12'hb27;
      20'h0f29c: out <= 12'hb27;
      20'h0f29d: out <= 12'hb27;
      20'h0f29e: out <= 12'hf87;
      20'h0f29f: out <= 12'hb27;
      20'h0f2a0: out <= 12'hee9;
      20'h0f2a1: out <= 12'hf87;
      20'h0f2a2: out <= 12'hee9;
      20'h0f2a3: out <= 12'hb27;
      20'h0f2a4: out <= 12'hb27;
      20'h0f2a5: out <= 12'hb27;
      20'h0f2a6: out <= 12'hf87;
      20'h0f2a7: out <= 12'hb27;
      20'h0f2a8: out <= 12'hee9;
      20'h0f2a9: out <= 12'hf87;
      20'h0f2aa: out <= 12'hee9;
      20'h0f2ab: out <= 12'hb27;
      20'h0f2ac: out <= 12'hb27;
      20'h0f2ad: out <= 12'hb27;
      20'h0f2ae: out <= 12'hf87;
      20'h0f2af: out <= 12'hb27;
      20'h0f2b0: out <= 12'hee9;
      20'h0f2b1: out <= 12'hf87;
      20'h0f2b2: out <= 12'hee9;
      20'h0f2b3: out <= 12'hb27;
      20'h0f2b4: out <= 12'hb27;
      20'h0f2b5: out <= 12'hb27;
      20'h0f2b6: out <= 12'hf87;
      20'h0f2b7: out <= 12'hb27;
      20'h0f2b8: out <= 12'hee9;
      20'h0f2b9: out <= 12'hf87;
      20'h0f2ba: out <= 12'hee9;
      20'h0f2bb: out <= 12'hb27;
      20'h0f2bc: out <= 12'hb27;
      20'h0f2bd: out <= 12'hb27;
      20'h0f2be: out <= 12'hf87;
      20'h0f2bf: out <= 12'hb27;
      20'h0f2c0: out <= 12'hee9;
      20'h0f2c1: out <= 12'hf87;
      20'h0f2c2: out <= 12'hee9;
      20'h0f2c3: out <= 12'hb27;
      20'h0f2c4: out <= 12'hb27;
      20'h0f2c5: out <= 12'hb27;
      20'h0f2c6: out <= 12'hf87;
      20'h0f2c7: out <= 12'hb27;
      20'h0f2c8: out <= 12'hee9;
      20'h0f2c9: out <= 12'hf87;
      20'h0f2ca: out <= 12'hee9;
      20'h0f2cb: out <= 12'hb27;
      20'h0f2cc: out <= 12'hb27;
      20'h0f2cd: out <= 12'hb27;
      20'h0f2ce: out <= 12'hf87;
      20'h0f2cf: out <= 12'hb27;
      20'h0f2d0: out <= 12'hfff;
      20'h0f2d1: out <= 12'hfff;
      20'h0f2d2: out <= 12'h666;
      20'h0f2d3: out <= 12'h666;
      20'h0f2d4: out <= 12'h666;
      20'h0f2d5: out <= 12'h666;
      20'h0f2d6: out <= 12'h666;
      20'h0f2d7: out <= 12'h666;
      20'h0f2d8: out <= 12'h666;
      20'h0f2d9: out <= 12'h666;
      20'h0f2da: out <= 12'h666;
      20'h0f2db: out <= 12'h666;
      20'h0f2dc: out <= 12'h666;
      20'h0f2dd: out <= 12'h666;
      20'h0f2de: out <= 12'h666;
      20'h0f2df: out <= 12'h666;
      20'h0f2e0: out <= 12'h666;
      20'h0f2e1: out <= 12'h666;
      20'h0f2e2: out <= 12'h666;
      20'h0f2e3: out <= 12'h666;
      20'h0f2e4: out <= 12'h666;
      20'h0f2e5: out <= 12'h666;
      20'h0f2e6: out <= 12'h666;
      20'h0f2e7: out <= 12'h666;
      20'h0f2e8: out <= 12'h666;
      20'h0f2e9: out <= 12'h666;
      20'h0f2ea: out <= 12'h666;
      20'h0f2eb: out <= 12'h666;
      20'h0f2ec: out <= 12'h666;
      20'h0f2ed: out <= 12'h666;
      20'h0f2ee: out <= 12'h666;
      20'h0f2ef: out <= 12'h666;
      20'h0f2f0: out <= 12'h666;
      20'h0f2f1: out <= 12'h666;
      20'h0f2f2: out <= 12'h666;
      20'h0f2f3: out <= 12'h666;
      20'h0f2f4: out <= 12'h666;
      20'h0f2f5: out <= 12'h666;
      20'h0f2f6: out <= 12'h666;
      20'h0f2f7: out <= 12'h666;
      20'h0f2f8: out <= 12'h666;
      20'h0f2f9: out <= 12'h666;
      20'h0f2fa: out <= 12'h666;
      20'h0f2fb: out <= 12'h666;
      20'h0f2fc: out <= 12'h666;
      20'h0f2fd: out <= 12'h666;
      20'h0f2fe: out <= 12'h666;
      20'h0f2ff: out <= 12'h666;
      20'h0f300: out <= 12'h603;
      20'h0f301: out <= 12'h603;
      20'h0f302: out <= 12'h603;
      20'h0f303: out <= 12'h603;
      20'h0f304: out <= 12'h603;
      20'h0f305: out <= 12'h603;
      20'h0f306: out <= 12'h603;
      20'h0f307: out <= 12'h603;
      20'h0f308: out <= 12'h603;
      20'h0f309: out <= 12'h603;
      20'h0f30a: out <= 12'h603;
      20'h0f30b: out <= 12'h603;
      20'h0f30c: out <= 12'h603;
      20'h0f30d: out <= 12'h603;
      20'h0f30e: out <= 12'h603;
      20'h0f30f: out <= 12'h603;
      20'h0f310: out <= 12'h603;
      20'h0f311: out <= 12'h603;
      20'h0f312: out <= 12'h603;
      20'h0f313: out <= 12'h603;
      20'h0f314: out <= 12'h603;
      20'h0f315: out <= 12'h603;
      20'h0f316: out <= 12'h603;
      20'h0f317: out <= 12'h603;
      20'h0f318: out <= 12'h603;
      20'h0f319: out <= 12'h603;
      20'h0f31a: out <= 12'h603;
      20'h0f31b: out <= 12'h603;
      20'h0f31c: out <= 12'h603;
      20'h0f31d: out <= 12'h603;
      20'h0f31e: out <= 12'h603;
      20'h0f31f: out <= 12'h603;
      20'h0f320: out <= 12'h603;
      20'h0f321: out <= 12'h603;
      20'h0f322: out <= 12'h603;
      20'h0f323: out <= 12'h603;
      20'h0f324: out <= 12'h603;
      20'h0f325: out <= 12'h603;
      20'h0f326: out <= 12'h603;
      20'h0f327: out <= 12'h603;
      20'h0f328: out <= 12'hfff;
      20'h0f329: out <= 12'hfff;
      20'h0f32a: out <= 12'h72f;
      20'h0f32b: out <= 12'h72f;
      20'h0f32c: out <= 12'h72f;
      20'h0f32d: out <= 12'h72f;
      20'h0f32e: out <= 12'h72f;
      20'h0f32f: out <= 12'h72f;
      20'h0f330: out <= 12'h72f;
      20'h0f331: out <= 12'h72f;
      20'h0f332: out <= 12'h72f;
      20'h0f333: out <= 12'h72f;
      20'h0f334: out <= 12'h72f;
      20'h0f335: out <= 12'h72f;
      20'h0f336: out <= 12'h72f;
      20'h0f337: out <= 12'h72f;
      20'h0f338: out <= 12'h72f;
      20'h0f339: out <= 12'h72f;
      20'h0f33a: out <= 12'h72f;
      20'h0f33b: out <= 12'h72f;
      20'h0f33c: out <= 12'h72f;
      20'h0f33d: out <= 12'h72f;
      20'h0f33e: out <= 12'h72f;
      20'h0f33f: out <= 12'h72f;
      20'h0f340: out <= 12'h72f;
      20'h0f341: out <= 12'h72f;
      20'h0f342: out <= 12'h72f;
      20'h0f343: out <= 12'h72f;
      20'h0f344: out <= 12'h72f;
      20'h0f345: out <= 12'h72f;
      20'h0f346: out <= 12'h72f;
      20'h0f347: out <= 12'h72f;
      20'h0f348: out <= 12'h72f;
      20'h0f349: out <= 12'h72f;
      20'h0f34a: out <= 12'h72f;
      20'h0f34b: out <= 12'h72f;
      20'h0f34c: out <= 12'h72f;
      20'h0f34d: out <= 12'h72f;
      20'h0f34e: out <= 12'h72f;
      20'h0f34f: out <= 12'h72f;
      20'h0f350: out <= 12'h603;
      20'h0f351: out <= 12'h603;
      20'h0f352: out <= 12'h603;
      20'h0f353: out <= 12'h603;
      20'h0f354: out <= 12'h603;
      20'h0f355: out <= 12'h603;
      20'h0f356: out <= 12'h603;
      20'h0f357: out <= 12'h603;
      20'h0f358: out <= 12'h603;
      20'h0f359: out <= 12'h603;
      20'h0f35a: out <= 12'h603;
      20'h0f35b: out <= 12'h603;
      20'h0f35c: out <= 12'h603;
      20'h0f35d: out <= 12'h603;
      20'h0f35e: out <= 12'h603;
      20'h0f35f: out <= 12'h603;
      20'h0f360: out <= 12'h603;
      20'h0f361: out <= 12'h603;
      20'h0f362: out <= 12'h603;
      20'h0f363: out <= 12'h603;
      20'h0f364: out <= 12'h603;
      20'h0f365: out <= 12'h603;
      20'h0f366: out <= 12'h603;
      20'h0f367: out <= 12'h603;
      20'h0f368: out <= 12'h603;
      20'h0f369: out <= 12'h603;
      20'h0f36a: out <= 12'h603;
      20'h0f36b: out <= 12'h603;
      20'h0f36c: out <= 12'h603;
      20'h0f36d: out <= 12'h603;
      20'h0f36e: out <= 12'h603;
      20'h0f36f: out <= 12'h603;
      20'h0f370: out <= 12'h603;
      20'h0f371: out <= 12'h603;
      20'h0f372: out <= 12'h603;
      20'h0f373: out <= 12'h603;
      20'h0f374: out <= 12'h603;
      20'h0f375: out <= 12'h603;
      20'h0f376: out <= 12'h603;
      20'h0f377: out <= 12'h603;
      20'h0f378: out <= 12'h603;
      20'h0f379: out <= 12'h603;
      20'h0f37a: out <= 12'h603;
      20'h0f37b: out <= 12'h603;
      20'h0f37c: out <= 12'h603;
      20'h0f37d: out <= 12'h603;
      20'h0f37e: out <= 12'h603;
      20'h0f37f: out <= 12'h603;
      20'h0f380: out <= 12'h603;
      20'h0f381: out <= 12'h603;
      20'h0f382: out <= 12'h603;
      20'h0f383: out <= 12'h603;
      20'h0f384: out <= 12'h603;
      20'h0f385: out <= 12'h603;
      20'h0f386: out <= 12'h603;
      20'h0f387: out <= 12'h603;
      20'h0f388: out <= 12'h603;
      20'h0f389: out <= 12'h603;
      20'h0f38a: out <= 12'h603;
      20'h0f38b: out <= 12'h603;
      20'h0f38c: out <= 12'h603;
      20'h0f38d: out <= 12'h603;
      20'h0f38e: out <= 12'h603;
      20'h0f38f: out <= 12'h603;
      20'h0f390: out <= 12'h603;
      20'h0f391: out <= 12'h603;
      20'h0f392: out <= 12'h603;
      20'h0f393: out <= 12'h603;
      20'h0f394: out <= 12'h603;
      20'h0f395: out <= 12'h603;
      20'h0f396: out <= 12'h603;
      20'h0f397: out <= 12'h603;
      20'h0f398: out <= 12'h603;
      20'h0f399: out <= 12'h603;
      20'h0f39a: out <= 12'h603;
      20'h0f39b: out <= 12'h603;
      20'h0f39c: out <= 12'h603;
      20'h0f39d: out <= 12'h603;
      20'h0f39e: out <= 12'h603;
      20'h0f39f: out <= 12'h603;
      20'h0f3a0: out <= 12'h603;
      20'h0f3a1: out <= 12'h603;
      20'h0f3a2: out <= 12'h603;
      20'h0f3a3: out <= 12'h603;
      20'h0f3a4: out <= 12'h603;
      20'h0f3a5: out <= 12'h603;
      20'h0f3a6: out <= 12'h603;
      20'h0f3a7: out <= 12'h603;
      20'h0f3a8: out <= 12'hee9;
      20'h0f3a9: out <= 12'hf87;
      20'h0f3aa: out <= 12'hf87;
      20'h0f3ab: out <= 12'hf87;
      20'h0f3ac: out <= 12'hf87;
      20'h0f3ad: out <= 12'hf87;
      20'h0f3ae: out <= 12'hf87;
      20'h0f3af: out <= 12'hb27;
      20'h0f3b0: out <= 12'hee9;
      20'h0f3b1: out <= 12'hf87;
      20'h0f3b2: out <= 12'hf87;
      20'h0f3b3: out <= 12'hf87;
      20'h0f3b4: out <= 12'hf87;
      20'h0f3b5: out <= 12'hf87;
      20'h0f3b6: out <= 12'hf87;
      20'h0f3b7: out <= 12'hb27;
      20'h0f3b8: out <= 12'hee9;
      20'h0f3b9: out <= 12'hf87;
      20'h0f3ba: out <= 12'hf87;
      20'h0f3bb: out <= 12'hf87;
      20'h0f3bc: out <= 12'hf87;
      20'h0f3bd: out <= 12'hf87;
      20'h0f3be: out <= 12'hf87;
      20'h0f3bf: out <= 12'hb27;
      20'h0f3c0: out <= 12'hee9;
      20'h0f3c1: out <= 12'hf87;
      20'h0f3c2: out <= 12'hf87;
      20'h0f3c3: out <= 12'hf87;
      20'h0f3c4: out <= 12'hf87;
      20'h0f3c5: out <= 12'hf87;
      20'h0f3c6: out <= 12'hf87;
      20'h0f3c7: out <= 12'hb27;
      20'h0f3c8: out <= 12'hee9;
      20'h0f3c9: out <= 12'hf87;
      20'h0f3ca: out <= 12'hf87;
      20'h0f3cb: out <= 12'hf87;
      20'h0f3cc: out <= 12'hf87;
      20'h0f3cd: out <= 12'hf87;
      20'h0f3ce: out <= 12'hf87;
      20'h0f3cf: out <= 12'hb27;
      20'h0f3d0: out <= 12'hee9;
      20'h0f3d1: out <= 12'hf87;
      20'h0f3d2: out <= 12'hf87;
      20'h0f3d3: out <= 12'hf87;
      20'h0f3d4: out <= 12'hf87;
      20'h0f3d5: out <= 12'hf87;
      20'h0f3d6: out <= 12'hf87;
      20'h0f3d7: out <= 12'hb27;
      20'h0f3d8: out <= 12'hee9;
      20'h0f3d9: out <= 12'hf87;
      20'h0f3da: out <= 12'hf87;
      20'h0f3db: out <= 12'hf87;
      20'h0f3dc: out <= 12'hf87;
      20'h0f3dd: out <= 12'hf87;
      20'h0f3de: out <= 12'hf87;
      20'h0f3df: out <= 12'hb27;
      20'h0f3e0: out <= 12'hee9;
      20'h0f3e1: out <= 12'hf87;
      20'h0f3e2: out <= 12'hf87;
      20'h0f3e3: out <= 12'hf87;
      20'h0f3e4: out <= 12'hf87;
      20'h0f3e5: out <= 12'hf87;
      20'h0f3e6: out <= 12'hf87;
      20'h0f3e7: out <= 12'hb27;
      20'h0f3e8: out <= 12'hfff;
      20'h0f3e9: out <= 12'h666;
      20'h0f3ea: out <= 12'h666;
      20'h0f3eb: out <= 12'h666;
      20'h0f3ec: out <= 12'h666;
      20'h0f3ed: out <= 12'h666;
      20'h0f3ee: out <= 12'h666;
      20'h0f3ef: out <= 12'h666;
      20'h0f3f0: out <= 12'h666;
      20'h0f3f1: out <= 12'h666;
      20'h0f3f2: out <= 12'h666;
      20'h0f3f3: out <= 12'h666;
      20'h0f3f4: out <= 12'h666;
      20'h0f3f5: out <= 12'h666;
      20'h0f3f6: out <= 12'h666;
      20'h0f3f7: out <= 12'h666;
      20'h0f3f8: out <= 12'h666;
      20'h0f3f9: out <= 12'h666;
      20'h0f3fa: out <= 12'h666;
      20'h0f3fb: out <= 12'h666;
      20'h0f3fc: out <= 12'h666;
      20'h0f3fd: out <= 12'h666;
      20'h0f3fe: out <= 12'h666;
      20'h0f3ff: out <= 12'h666;
      20'h0f400: out <= 12'h666;
      20'h0f401: out <= 12'h666;
      20'h0f402: out <= 12'h666;
      20'h0f403: out <= 12'h666;
      20'h0f404: out <= 12'h666;
      20'h0f405: out <= 12'h666;
      20'h0f406: out <= 12'h666;
      20'h0f407: out <= 12'h666;
      20'h0f408: out <= 12'h666;
      20'h0f409: out <= 12'h666;
      20'h0f40a: out <= 12'h666;
      20'h0f40b: out <= 12'h666;
      20'h0f40c: out <= 12'h666;
      20'h0f40d: out <= 12'h666;
      20'h0f40e: out <= 12'h666;
      20'h0f40f: out <= 12'h666;
      20'h0f410: out <= 12'h666;
      20'h0f411: out <= 12'h666;
      20'h0f412: out <= 12'h666;
      20'h0f413: out <= 12'h666;
      20'h0f414: out <= 12'h666;
      20'h0f415: out <= 12'h666;
      20'h0f416: out <= 12'h666;
      20'h0f417: out <= 12'h666;
      20'h0f418: out <= 12'h603;
      20'h0f419: out <= 12'h603;
      20'h0f41a: out <= 12'h603;
      20'h0f41b: out <= 12'h603;
      20'h0f41c: out <= 12'h603;
      20'h0f41d: out <= 12'h603;
      20'h0f41e: out <= 12'h603;
      20'h0f41f: out <= 12'h603;
      20'h0f420: out <= 12'h603;
      20'h0f421: out <= 12'h603;
      20'h0f422: out <= 12'h603;
      20'h0f423: out <= 12'h603;
      20'h0f424: out <= 12'h603;
      20'h0f425: out <= 12'h603;
      20'h0f426: out <= 12'h603;
      20'h0f427: out <= 12'h603;
      20'h0f428: out <= 12'h603;
      20'h0f429: out <= 12'h603;
      20'h0f42a: out <= 12'h603;
      20'h0f42b: out <= 12'h603;
      20'h0f42c: out <= 12'h603;
      20'h0f42d: out <= 12'h603;
      20'h0f42e: out <= 12'h603;
      20'h0f42f: out <= 12'h603;
      20'h0f430: out <= 12'h603;
      20'h0f431: out <= 12'h603;
      20'h0f432: out <= 12'h603;
      20'h0f433: out <= 12'h603;
      20'h0f434: out <= 12'h603;
      20'h0f435: out <= 12'h603;
      20'h0f436: out <= 12'h603;
      20'h0f437: out <= 12'h603;
      20'h0f438: out <= 12'h603;
      20'h0f439: out <= 12'h603;
      20'h0f43a: out <= 12'h603;
      20'h0f43b: out <= 12'h603;
      20'h0f43c: out <= 12'h603;
      20'h0f43d: out <= 12'h603;
      20'h0f43e: out <= 12'h603;
      20'h0f43f: out <= 12'h603;
      20'h0f440: out <= 12'hfff;
      20'h0f441: out <= 12'h72f;
      20'h0f442: out <= 12'h72f;
      20'h0f443: out <= 12'h72f;
      20'h0f444: out <= 12'h72f;
      20'h0f445: out <= 12'h72f;
      20'h0f446: out <= 12'h72f;
      20'h0f447: out <= 12'h72f;
      20'h0f448: out <= 12'h72f;
      20'h0f449: out <= 12'h72f;
      20'h0f44a: out <= 12'h72f;
      20'h0f44b: out <= 12'h72f;
      20'h0f44c: out <= 12'h72f;
      20'h0f44d: out <= 12'h72f;
      20'h0f44e: out <= 12'h72f;
      20'h0f44f: out <= 12'h72f;
      20'h0f450: out <= 12'h72f;
      20'h0f451: out <= 12'h72f;
      20'h0f452: out <= 12'h72f;
      20'h0f453: out <= 12'h72f;
      20'h0f454: out <= 12'h72f;
      20'h0f455: out <= 12'h72f;
      20'h0f456: out <= 12'h72f;
      20'h0f457: out <= 12'h72f;
      20'h0f458: out <= 12'h72f;
      20'h0f459: out <= 12'h72f;
      20'h0f45a: out <= 12'h72f;
      20'h0f45b: out <= 12'h72f;
      20'h0f45c: out <= 12'h72f;
      20'h0f45d: out <= 12'h72f;
      20'h0f45e: out <= 12'h72f;
      20'h0f45f: out <= 12'h72f;
      20'h0f460: out <= 12'h72f;
      20'h0f461: out <= 12'h72f;
      20'h0f462: out <= 12'h72f;
      20'h0f463: out <= 12'h72f;
      20'h0f464: out <= 12'h72f;
      20'h0f465: out <= 12'h72f;
      20'h0f466: out <= 12'h72f;
      20'h0f467: out <= 12'h72f;
      20'h0f468: out <= 12'h603;
      20'h0f469: out <= 12'h603;
      20'h0f46a: out <= 12'h603;
      20'h0f46b: out <= 12'h603;
      20'h0f46c: out <= 12'h603;
      20'h0f46d: out <= 12'h603;
      20'h0f46e: out <= 12'h603;
      20'h0f46f: out <= 12'h603;
      20'h0f470: out <= 12'h603;
      20'h0f471: out <= 12'h603;
      20'h0f472: out <= 12'h603;
      20'h0f473: out <= 12'h603;
      20'h0f474: out <= 12'h603;
      20'h0f475: out <= 12'h603;
      20'h0f476: out <= 12'h603;
      20'h0f477: out <= 12'h603;
      20'h0f478: out <= 12'h603;
      20'h0f479: out <= 12'h603;
      20'h0f47a: out <= 12'h603;
      20'h0f47b: out <= 12'h603;
      20'h0f47c: out <= 12'h603;
      20'h0f47d: out <= 12'h603;
      20'h0f47e: out <= 12'h603;
      20'h0f47f: out <= 12'h603;
      20'h0f480: out <= 12'h603;
      20'h0f481: out <= 12'h603;
      20'h0f482: out <= 12'h603;
      20'h0f483: out <= 12'h603;
      20'h0f484: out <= 12'h603;
      20'h0f485: out <= 12'h603;
      20'h0f486: out <= 12'h603;
      20'h0f487: out <= 12'h603;
      20'h0f488: out <= 12'h603;
      20'h0f489: out <= 12'h603;
      20'h0f48a: out <= 12'h603;
      20'h0f48b: out <= 12'h603;
      20'h0f48c: out <= 12'h603;
      20'h0f48d: out <= 12'h603;
      20'h0f48e: out <= 12'h603;
      20'h0f48f: out <= 12'h603;
      20'h0f490: out <= 12'h603;
      20'h0f491: out <= 12'h603;
      20'h0f492: out <= 12'h603;
      20'h0f493: out <= 12'h603;
      20'h0f494: out <= 12'h603;
      20'h0f495: out <= 12'h603;
      20'h0f496: out <= 12'h603;
      20'h0f497: out <= 12'h603;
      20'h0f498: out <= 12'h603;
      20'h0f499: out <= 12'h603;
      20'h0f49a: out <= 12'h603;
      20'h0f49b: out <= 12'h603;
      20'h0f49c: out <= 12'h603;
      20'h0f49d: out <= 12'h603;
      20'h0f49e: out <= 12'h603;
      20'h0f49f: out <= 12'h603;
      20'h0f4a0: out <= 12'h603;
      20'h0f4a1: out <= 12'h603;
      20'h0f4a2: out <= 12'h603;
      20'h0f4a3: out <= 12'h603;
      20'h0f4a4: out <= 12'h603;
      20'h0f4a5: out <= 12'h603;
      20'h0f4a6: out <= 12'h603;
      20'h0f4a7: out <= 12'h603;
      20'h0f4a8: out <= 12'h603;
      20'h0f4a9: out <= 12'h603;
      20'h0f4aa: out <= 12'h603;
      20'h0f4ab: out <= 12'h603;
      20'h0f4ac: out <= 12'h603;
      20'h0f4ad: out <= 12'h603;
      20'h0f4ae: out <= 12'h603;
      20'h0f4af: out <= 12'h603;
      20'h0f4b0: out <= 12'h603;
      20'h0f4b1: out <= 12'h603;
      20'h0f4b2: out <= 12'h603;
      20'h0f4b3: out <= 12'h603;
      20'h0f4b4: out <= 12'h603;
      20'h0f4b5: out <= 12'h603;
      20'h0f4b6: out <= 12'h603;
      20'h0f4b7: out <= 12'h603;
      20'h0f4b8: out <= 12'h603;
      20'h0f4b9: out <= 12'h